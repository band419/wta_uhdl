//[UHDL]Content Start [md5:6e927582602471e237b52f7140ea2183]
module WtaTree_num_pp_10_pp_width_32 (
	input  [31:0] pp_0,
	input  [31:0] pp_1,
	input  [31:0] pp_2,
	input  [31:0] pp_3,
	input  [31:0] pp_4,
	input  [31:0] pp_5,
	input  [31:0] pp_6,
	input  [31:0] pp_7,
	input  [31:0] pp_8,
	input  [31:0] pp_9,
	output [31:0] ps_0,
	output [31:0] ps_1);

	//Wire define for this module.
	wire [0:0] p_0_0                ;
	wire [0:0] p_0_1                ;
	wire [0:0] p_0_2                ;
	wire [0:0] p_0_3                ;
	wire [0:0] p_0_4                ;
	wire [0:0] p_0_5                ;
	wire [0:0] p_0_6                ;
	wire [0:0] p_0_7                ;
	wire [0:0] p_0_8                ;
	wire [0:0] p_0_9                ;
	wire [0:0] p_0_10               ;
	wire [0:0] p_0_11               ;
	wire [0:0] p_0_12               ;
	wire [0:0] p_0_13               ;
	wire [0:0] p_0_14               ;
	wire [0:0] p_0_15               ;
	wire [0:0] p_0_16               ;
	wire [0:0] p_0_17               ;
	wire [0:0] p_0_18               ;
	wire [0:0] p_0_19               ;
	wire [0:0] p_0_20               ;
	wire [0:0] p_0_21               ;
	wire [0:0] p_0_22               ;
	wire [0:0] p_0_23               ;
	wire [0:0] p_0_24               ;
	wire [0:0] p_0_25               ;
	wire [0:0] p_0_26               ;
	wire [0:0] p_0_27               ;
	wire [0:0] p_0_28               ;
	wire [0:0] p_0_29               ;
	wire [0:0] p_0_30               ;
	wire [0:0] p_0_31               ;
	wire [0:0] p_1_0                ;
	wire [0:0] p_1_1                ;
	wire [0:0] p_1_2                ;
	wire [0:0] p_1_3                ;
	wire [0:0] p_1_4                ;
	wire [0:0] p_1_5                ;
	wire [0:0] p_1_6                ;
	wire [0:0] p_1_7                ;
	wire [0:0] p_1_8                ;
	wire [0:0] p_1_9                ;
	wire [0:0] p_1_10               ;
	wire [0:0] p_1_11               ;
	wire [0:0] p_1_12               ;
	wire [0:0] p_1_13               ;
	wire [0:0] p_1_14               ;
	wire [0:0] p_1_15               ;
	wire [0:0] p_1_16               ;
	wire [0:0] p_1_17               ;
	wire [0:0] p_1_18               ;
	wire [0:0] p_1_19               ;
	wire [0:0] p_1_20               ;
	wire [0:0] p_1_21               ;
	wire [0:0] p_1_22               ;
	wire [0:0] p_1_23               ;
	wire [0:0] p_1_24               ;
	wire [0:0] p_1_25               ;
	wire [0:0] p_1_26               ;
	wire [0:0] p_1_27               ;
	wire [0:0] p_1_28               ;
	wire [0:0] p_1_29               ;
	wire [0:0] p_1_30               ;
	wire [0:0] p_1_31               ;
	wire [0:0] p_2_0                ;
	wire [0:0] p_2_1                ;
	wire [0:0] p_2_2                ;
	wire [0:0] p_2_3                ;
	wire [0:0] p_2_4                ;
	wire [0:0] p_2_5                ;
	wire [0:0] p_2_6                ;
	wire [0:0] p_2_7                ;
	wire [0:0] p_2_8                ;
	wire [0:0] p_2_9                ;
	wire [0:0] p_2_10               ;
	wire [0:0] p_2_11               ;
	wire [0:0] p_2_12               ;
	wire [0:0] p_2_13               ;
	wire [0:0] p_2_14               ;
	wire [0:0] p_2_15               ;
	wire [0:0] p_2_16               ;
	wire [0:0] p_2_17               ;
	wire [0:0] p_2_18               ;
	wire [0:0] p_2_19               ;
	wire [0:0] p_2_20               ;
	wire [0:0] p_2_21               ;
	wire [0:0] p_2_22               ;
	wire [0:0] p_2_23               ;
	wire [0:0] p_2_24               ;
	wire [0:0] p_2_25               ;
	wire [0:0] p_2_26               ;
	wire [0:0] p_2_27               ;
	wire [0:0] p_2_28               ;
	wire [0:0] p_2_29               ;
	wire [0:0] p_2_30               ;
	wire [0:0] p_2_31               ;
	wire [0:0] p_3_0                ;
	wire [0:0] p_3_1                ;
	wire [0:0] p_3_2                ;
	wire [0:0] p_3_3                ;
	wire [0:0] p_3_4                ;
	wire [0:0] p_3_5                ;
	wire [0:0] p_3_6                ;
	wire [0:0] p_3_7                ;
	wire [0:0] p_3_8                ;
	wire [0:0] p_3_9                ;
	wire [0:0] p_3_10               ;
	wire [0:0] p_3_11               ;
	wire [0:0] p_3_12               ;
	wire [0:0] p_3_13               ;
	wire [0:0] p_3_14               ;
	wire [0:0] p_3_15               ;
	wire [0:0] p_3_16               ;
	wire [0:0] p_3_17               ;
	wire [0:0] p_3_18               ;
	wire [0:0] p_3_19               ;
	wire [0:0] p_3_20               ;
	wire [0:0] p_3_21               ;
	wire [0:0] p_3_22               ;
	wire [0:0] p_3_23               ;
	wire [0:0] p_3_24               ;
	wire [0:0] p_3_25               ;
	wire [0:0] p_3_26               ;
	wire [0:0] p_3_27               ;
	wire [0:0] p_3_28               ;
	wire [0:0] p_3_29               ;
	wire [0:0] p_3_30               ;
	wire [0:0] p_3_31               ;
	wire [0:0] p_4_0                ;
	wire [0:0] p_4_1                ;
	wire [0:0] p_4_2                ;
	wire [0:0] p_4_3                ;
	wire [0:0] p_4_4                ;
	wire [0:0] p_4_5                ;
	wire [0:0] p_4_6                ;
	wire [0:0] p_4_7                ;
	wire [0:0] p_4_8                ;
	wire [0:0] p_4_9                ;
	wire [0:0] p_4_10               ;
	wire [0:0] p_4_11               ;
	wire [0:0] p_4_12               ;
	wire [0:0] p_4_13               ;
	wire [0:0] p_4_14               ;
	wire [0:0] p_4_15               ;
	wire [0:0] p_4_16               ;
	wire [0:0] p_4_17               ;
	wire [0:0] p_4_18               ;
	wire [0:0] p_4_19               ;
	wire [0:0] p_4_20               ;
	wire [0:0] p_4_21               ;
	wire [0:0] p_4_22               ;
	wire [0:0] p_4_23               ;
	wire [0:0] p_4_24               ;
	wire [0:0] p_4_25               ;
	wire [0:0] p_4_26               ;
	wire [0:0] p_4_27               ;
	wire [0:0] p_4_28               ;
	wire [0:0] p_4_29               ;
	wire [0:0] p_4_30               ;
	wire [0:0] p_4_31               ;
	wire [0:0] p_5_0                ;
	wire [0:0] p_5_1                ;
	wire [0:0] p_5_2                ;
	wire [0:0] p_5_3                ;
	wire [0:0] p_5_4                ;
	wire [0:0] p_5_5                ;
	wire [0:0] p_5_6                ;
	wire [0:0] p_5_7                ;
	wire [0:0] p_5_8                ;
	wire [0:0] p_5_9                ;
	wire [0:0] p_5_10               ;
	wire [0:0] p_5_11               ;
	wire [0:0] p_5_12               ;
	wire [0:0] p_5_13               ;
	wire [0:0] p_5_14               ;
	wire [0:0] p_5_15               ;
	wire [0:0] p_5_16               ;
	wire [0:0] p_5_17               ;
	wire [0:0] p_5_18               ;
	wire [0:0] p_5_19               ;
	wire [0:0] p_5_20               ;
	wire [0:0] p_5_21               ;
	wire [0:0] p_5_22               ;
	wire [0:0] p_5_23               ;
	wire [0:0] p_5_24               ;
	wire [0:0] p_5_25               ;
	wire [0:0] p_5_26               ;
	wire [0:0] p_5_27               ;
	wire [0:0] p_5_28               ;
	wire [0:0] p_5_29               ;
	wire [0:0] p_5_30               ;
	wire [0:0] p_5_31               ;
	wire [0:0] p_6_0                ;
	wire [0:0] p_6_1                ;
	wire [0:0] p_6_2                ;
	wire [0:0] p_6_3                ;
	wire [0:0] p_6_4                ;
	wire [0:0] p_6_5                ;
	wire [0:0] p_6_6                ;
	wire [0:0] p_6_7                ;
	wire [0:0] p_6_8                ;
	wire [0:0] p_6_9                ;
	wire [0:0] p_6_10               ;
	wire [0:0] p_6_11               ;
	wire [0:0] p_6_12               ;
	wire [0:0] p_6_13               ;
	wire [0:0] p_6_14               ;
	wire [0:0] p_6_15               ;
	wire [0:0] p_6_16               ;
	wire [0:0] p_6_17               ;
	wire [0:0] p_6_18               ;
	wire [0:0] p_6_19               ;
	wire [0:0] p_6_20               ;
	wire [0:0] p_6_21               ;
	wire [0:0] p_6_22               ;
	wire [0:0] p_6_23               ;
	wire [0:0] p_6_24               ;
	wire [0:0] p_6_25               ;
	wire [0:0] p_6_26               ;
	wire [0:0] p_6_27               ;
	wire [0:0] p_6_28               ;
	wire [0:0] p_6_29               ;
	wire [0:0] p_6_30               ;
	wire [0:0] p_6_31               ;
	wire [0:0] p_7_0                ;
	wire [0:0] p_7_1                ;
	wire [0:0] p_7_2                ;
	wire [0:0] p_7_3                ;
	wire [0:0] p_7_4                ;
	wire [0:0] p_7_5                ;
	wire [0:0] p_7_6                ;
	wire [0:0] p_7_7                ;
	wire [0:0] p_7_8                ;
	wire [0:0] p_7_9                ;
	wire [0:0] p_7_10               ;
	wire [0:0] p_7_11               ;
	wire [0:0] p_7_12               ;
	wire [0:0] p_7_13               ;
	wire [0:0] p_7_14               ;
	wire [0:0] p_7_15               ;
	wire [0:0] p_7_16               ;
	wire [0:0] p_7_17               ;
	wire [0:0] p_7_18               ;
	wire [0:0] p_7_19               ;
	wire [0:0] p_7_20               ;
	wire [0:0] p_7_21               ;
	wire [0:0] p_7_22               ;
	wire [0:0] p_7_23               ;
	wire [0:0] p_7_24               ;
	wire [0:0] p_7_25               ;
	wire [0:0] p_7_26               ;
	wire [0:0] p_7_27               ;
	wire [0:0] p_7_28               ;
	wire [0:0] p_7_29               ;
	wire [0:0] p_7_30               ;
	wire [0:0] p_7_31               ;
	wire [0:0] p_8_0                ;
	wire [0:0] p_8_1                ;
	wire [0:0] p_8_2                ;
	wire [0:0] p_8_3                ;
	wire [0:0] p_8_4                ;
	wire [0:0] p_8_5                ;
	wire [0:0] p_8_6                ;
	wire [0:0] p_8_7                ;
	wire [0:0] p_8_8                ;
	wire [0:0] p_8_9                ;
	wire [0:0] p_8_10               ;
	wire [0:0] p_8_11               ;
	wire [0:0] p_8_12               ;
	wire [0:0] p_8_13               ;
	wire [0:0] p_8_14               ;
	wire [0:0] p_8_15               ;
	wire [0:0] p_8_16               ;
	wire [0:0] p_8_17               ;
	wire [0:0] p_8_18               ;
	wire [0:0] p_8_19               ;
	wire [0:0] p_8_20               ;
	wire [0:0] p_8_21               ;
	wire [0:0] p_8_22               ;
	wire [0:0] p_8_23               ;
	wire [0:0] p_8_24               ;
	wire [0:0] p_8_25               ;
	wire [0:0] p_8_26               ;
	wire [0:0] p_8_27               ;
	wire [0:0] p_8_28               ;
	wire [0:0] p_8_29               ;
	wire [0:0] p_8_30               ;
	wire [0:0] p_8_31               ;
	wire [0:0] p_9_0                ;
	wire [0:0] p_9_1                ;
	wire [0:0] p_9_2                ;
	wire [0:0] p_9_3                ;
	wire [0:0] p_9_4                ;
	wire [0:0] p_9_5                ;
	wire [0:0] p_9_6                ;
	wire [0:0] p_9_7                ;
	wire [0:0] p_9_8                ;
	wire [0:0] p_9_9                ;
	wire [0:0] p_9_10               ;
	wire [0:0] p_9_11               ;
	wire [0:0] p_9_12               ;
	wire [0:0] p_9_13               ;
	wire [0:0] p_9_14               ;
	wire [0:0] p_9_15               ;
	wire [0:0] p_9_16               ;
	wire [0:0] p_9_17               ;
	wire [0:0] p_9_18               ;
	wire [0:0] p_9_19               ;
	wire [0:0] p_9_20               ;
	wire [0:0] p_9_21               ;
	wire [0:0] p_9_22               ;
	wire [0:0] p_9_23               ;
	wire [0:0] p_9_24               ;
	wire [0:0] p_9_25               ;
	wire [0:0] p_9_26               ;
	wire [0:0] p_9_27               ;
	wire [0:0] p_9_28               ;
	wire [0:0] p_9_29               ;
	wire [0:0] p_9_30               ;
	wire [0:0] p_9_31               ;
	wire [0:0] comp_l0_p0_col0_cout ;
	wire [0:0] comp_l0_p0_col0_sum  ;
	wire [0:0] comp_l0_p0_col1_cout ;
	wire [0:0] comp_l0_p0_col1_sum  ;
	wire [0:0] comp_l0_p0_col2_cout ;
	wire [0:0] comp_l0_p0_col2_sum  ;
	wire [0:0] comp_l0_p0_col3_cout ;
	wire [0:0] comp_l0_p0_col3_sum  ;
	wire [0:0] comp_l0_p0_col4_cout ;
	wire [0:0] comp_l0_p0_col4_sum  ;
	wire [0:0] comp_l0_p0_col5_cout ;
	wire [0:0] comp_l0_p0_col5_sum  ;
	wire [0:0] comp_l0_p0_col6_cout ;
	wire [0:0] comp_l0_p0_col6_sum  ;
	wire [0:0] comp_l0_p0_col7_cout ;
	wire [0:0] comp_l0_p0_col7_sum  ;
	wire [0:0] comp_l0_p0_col8_cout ;
	wire [0:0] comp_l0_p0_col8_sum  ;
	wire [0:0] comp_l0_p0_col9_cout ;
	wire [0:0] comp_l0_p0_col9_sum  ;
	wire [0:0] comp_l0_p0_col10_cout;
	wire [0:0] comp_l0_p0_col10_sum ;
	wire [0:0] comp_l0_p0_col11_cout;
	wire [0:0] comp_l0_p0_col11_sum ;
	wire [0:0] comp_l0_p0_col12_cout;
	wire [0:0] comp_l0_p0_col12_sum ;
	wire [0:0] comp_l0_p0_col13_cout;
	wire [0:0] comp_l0_p0_col13_sum ;
	wire [0:0] comp_l0_p0_col14_cout;
	wire [0:0] comp_l0_p0_col14_sum ;
	wire [0:0] comp_l0_p0_col15_cout;
	wire [0:0] comp_l0_p0_col15_sum ;
	wire [0:0] comp_l0_p0_col16_cout;
	wire [0:0] comp_l0_p0_col16_sum ;
	wire [0:0] comp_l0_p0_col17_cout;
	wire [0:0] comp_l0_p0_col17_sum ;
	wire [0:0] comp_l0_p0_col18_cout;
	wire [0:0] comp_l0_p0_col18_sum ;
	wire [0:0] comp_l0_p0_col19_cout;
	wire [0:0] comp_l0_p0_col19_sum ;
	wire [0:0] comp_l0_p0_col20_cout;
	wire [0:0] comp_l0_p0_col20_sum ;
	wire [0:0] comp_l0_p0_col21_cout;
	wire [0:0] comp_l0_p0_col21_sum ;
	wire [0:0] comp_l0_p0_col22_cout;
	wire [0:0] comp_l0_p0_col22_sum ;
	wire [0:0] comp_l0_p0_col23_cout;
	wire [0:0] comp_l0_p0_col23_sum ;
	wire [0:0] comp_l0_p0_col24_cout;
	wire [0:0] comp_l0_p0_col24_sum ;
	wire [0:0] comp_l0_p0_col25_cout;
	wire [0:0] comp_l0_p0_col25_sum ;
	wire [0:0] comp_l0_p0_col26_cout;
	wire [0:0] comp_l0_p0_col26_sum ;
	wire [0:0] comp_l0_p0_col27_cout;
	wire [0:0] comp_l0_p0_col27_sum ;
	wire [0:0] comp_l0_p0_col28_cout;
	wire [0:0] comp_l0_p0_col28_sum ;
	wire [0:0] comp_l0_p0_col29_cout;
	wire [0:0] comp_l0_p0_col29_sum ;
	wire [0:0] comp_l0_p0_col30_cout;
	wire [0:0] comp_l0_p0_col30_sum ;
	wire [0:0] comp_l0_p0_col31_cout;
	wire [0:0] comp_l0_p0_col31_sum ;
	wire [0:0] comp_pad_l0_p0       ;
	wire [0:0] comp_l0_p1_col0_cout ;
	wire [0:0] comp_l0_p1_col0_sum  ;
	wire [0:0] comp_l0_p1_col1_cout ;
	wire [0:0] comp_l0_p1_col1_sum  ;
	wire [0:0] comp_l0_p1_col2_cout ;
	wire [0:0] comp_l0_p1_col2_sum  ;
	wire [0:0] comp_l0_p1_col3_cout ;
	wire [0:0] comp_l0_p1_col3_sum  ;
	wire [0:0] comp_l0_p1_col4_cout ;
	wire [0:0] comp_l0_p1_col4_sum  ;
	wire [0:0] comp_l0_p1_col5_cout ;
	wire [0:0] comp_l0_p1_col5_sum  ;
	wire [0:0] comp_l0_p1_col6_cout ;
	wire [0:0] comp_l0_p1_col6_sum  ;
	wire [0:0] comp_l0_p1_col7_cout ;
	wire [0:0] comp_l0_p1_col7_sum  ;
	wire [0:0] comp_l0_p1_col8_cout ;
	wire [0:0] comp_l0_p1_col8_sum  ;
	wire [0:0] comp_l0_p1_col9_cout ;
	wire [0:0] comp_l0_p1_col9_sum  ;
	wire [0:0] comp_l0_p1_col10_cout;
	wire [0:0] comp_l0_p1_col10_sum ;
	wire [0:0] comp_l0_p1_col11_cout;
	wire [0:0] comp_l0_p1_col11_sum ;
	wire [0:0] comp_l0_p1_col12_cout;
	wire [0:0] comp_l0_p1_col12_sum ;
	wire [0:0] comp_l0_p1_col13_cout;
	wire [0:0] comp_l0_p1_col13_sum ;
	wire [0:0] comp_l0_p1_col14_cout;
	wire [0:0] comp_l0_p1_col14_sum ;
	wire [0:0] comp_l0_p1_col15_cout;
	wire [0:0] comp_l0_p1_col15_sum ;
	wire [0:0] comp_l0_p1_col16_cout;
	wire [0:0] comp_l0_p1_col16_sum ;
	wire [0:0] comp_l0_p1_col17_cout;
	wire [0:0] comp_l0_p1_col17_sum ;
	wire [0:0] comp_l0_p1_col18_cout;
	wire [0:0] comp_l0_p1_col18_sum ;
	wire [0:0] comp_l0_p1_col19_cout;
	wire [0:0] comp_l0_p1_col19_sum ;
	wire [0:0] comp_l0_p1_col20_cout;
	wire [0:0] comp_l0_p1_col20_sum ;
	wire [0:0] comp_l0_p1_col21_cout;
	wire [0:0] comp_l0_p1_col21_sum ;
	wire [0:0] comp_l0_p1_col22_cout;
	wire [0:0] comp_l0_p1_col22_sum ;
	wire [0:0] comp_l0_p1_col23_cout;
	wire [0:0] comp_l0_p1_col23_sum ;
	wire [0:0] comp_l0_p1_col24_cout;
	wire [0:0] comp_l0_p1_col24_sum ;
	wire [0:0] comp_l0_p1_col25_cout;
	wire [0:0] comp_l0_p1_col25_sum ;
	wire [0:0] comp_l0_p1_col26_cout;
	wire [0:0] comp_l0_p1_col26_sum ;
	wire [0:0] comp_l0_p1_col27_cout;
	wire [0:0] comp_l0_p1_col27_sum ;
	wire [0:0] comp_l0_p1_col28_cout;
	wire [0:0] comp_l0_p1_col28_sum ;
	wire [0:0] comp_l0_p1_col29_cout;
	wire [0:0] comp_l0_p1_col29_sum ;
	wire [0:0] comp_l0_p1_col30_cout;
	wire [0:0] comp_l0_p1_col30_sum ;
	wire [0:0] comp_l0_p1_col31_cout;
	wire [0:0] comp_l0_p1_col31_sum ;
	wire [0:0] comp_pad_l0_p1       ;
	wire [0:0] comp_l0_p2_col0_cout ;
	wire [0:0] comp_l0_p2_col0_sum  ;
	wire [0:0] comp_l0_p2_col1_cout ;
	wire [0:0] comp_l0_p2_col1_sum  ;
	wire [0:0] comp_l0_p2_col2_cout ;
	wire [0:0] comp_l0_p2_col2_sum  ;
	wire [0:0] comp_l0_p2_col3_cout ;
	wire [0:0] comp_l0_p2_col3_sum  ;
	wire [0:0] comp_l0_p2_col4_cout ;
	wire [0:0] comp_l0_p2_col4_sum  ;
	wire [0:0] comp_l0_p2_col5_cout ;
	wire [0:0] comp_l0_p2_col5_sum  ;
	wire [0:0] comp_l0_p2_col6_cout ;
	wire [0:0] comp_l0_p2_col6_sum  ;
	wire [0:0] comp_l0_p2_col7_cout ;
	wire [0:0] comp_l0_p2_col7_sum  ;
	wire [0:0] comp_l0_p2_col8_cout ;
	wire [0:0] comp_l0_p2_col8_sum  ;
	wire [0:0] comp_l0_p2_col9_cout ;
	wire [0:0] comp_l0_p2_col9_sum  ;
	wire [0:0] comp_l0_p2_col10_cout;
	wire [0:0] comp_l0_p2_col10_sum ;
	wire [0:0] comp_l0_p2_col11_cout;
	wire [0:0] comp_l0_p2_col11_sum ;
	wire [0:0] comp_l0_p2_col12_cout;
	wire [0:0] comp_l0_p2_col12_sum ;
	wire [0:0] comp_l0_p2_col13_cout;
	wire [0:0] comp_l0_p2_col13_sum ;
	wire [0:0] comp_l0_p2_col14_cout;
	wire [0:0] comp_l0_p2_col14_sum ;
	wire [0:0] comp_l0_p2_col15_cout;
	wire [0:0] comp_l0_p2_col15_sum ;
	wire [0:0] comp_l0_p2_col16_cout;
	wire [0:0] comp_l0_p2_col16_sum ;
	wire [0:0] comp_l0_p2_col17_cout;
	wire [0:0] comp_l0_p2_col17_sum ;
	wire [0:0] comp_l0_p2_col18_cout;
	wire [0:0] comp_l0_p2_col18_sum ;
	wire [0:0] comp_l0_p2_col19_cout;
	wire [0:0] comp_l0_p2_col19_sum ;
	wire [0:0] comp_l0_p2_col20_cout;
	wire [0:0] comp_l0_p2_col20_sum ;
	wire [0:0] comp_l0_p2_col21_cout;
	wire [0:0] comp_l0_p2_col21_sum ;
	wire [0:0] comp_l0_p2_col22_cout;
	wire [0:0] comp_l0_p2_col22_sum ;
	wire [0:0] comp_l0_p2_col23_cout;
	wire [0:0] comp_l0_p2_col23_sum ;
	wire [0:0] comp_l0_p2_col24_cout;
	wire [0:0] comp_l0_p2_col24_sum ;
	wire [0:0] comp_l0_p2_col25_cout;
	wire [0:0] comp_l0_p2_col25_sum ;
	wire [0:0] comp_l0_p2_col26_cout;
	wire [0:0] comp_l0_p2_col26_sum ;
	wire [0:0] comp_l0_p2_col27_cout;
	wire [0:0] comp_l0_p2_col27_sum ;
	wire [0:0] comp_l0_p2_col28_cout;
	wire [0:0] comp_l0_p2_col28_sum ;
	wire [0:0] comp_l0_p2_col29_cout;
	wire [0:0] comp_l0_p2_col29_sum ;
	wire [0:0] comp_l0_p2_col30_cout;
	wire [0:0] comp_l0_p2_col30_sum ;
	wire [0:0] comp_l0_p2_col31_cout;
	wire [0:0] comp_l0_p2_col31_sum ;
	wire [0:0] comp_pad_l0_p2       ;
	wire [0:0] comp_l1_p0_col0_cout ;
	wire [0:0] comp_l1_p0_col0_sum  ;
	wire [0:0] comp_l1_p0_col1_cout ;
	wire [0:0] comp_l1_p0_col1_sum  ;
	wire [0:0] comp_l1_p0_col2_cout ;
	wire [0:0] comp_l1_p0_col2_sum  ;
	wire [0:0] comp_l1_p0_col3_cout ;
	wire [0:0] comp_l1_p0_col3_sum  ;
	wire [0:0] comp_l1_p0_col4_cout ;
	wire [0:0] comp_l1_p0_col4_sum  ;
	wire [0:0] comp_l1_p0_col5_cout ;
	wire [0:0] comp_l1_p0_col5_sum  ;
	wire [0:0] comp_l1_p0_col6_cout ;
	wire [0:0] comp_l1_p0_col6_sum  ;
	wire [0:0] comp_l1_p0_col7_cout ;
	wire [0:0] comp_l1_p0_col7_sum  ;
	wire [0:0] comp_l1_p0_col8_cout ;
	wire [0:0] comp_l1_p0_col8_sum  ;
	wire [0:0] comp_l1_p0_col9_cout ;
	wire [0:0] comp_l1_p0_col9_sum  ;
	wire [0:0] comp_l1_p0_col10_cout;
	wire [0:0] comp_l1_p0_col10_sum ;
	wire [0:0] comp_l1_p0_col11_cout;
	wire [0:0] comp_l1_p0_col11_sum ;
	wire [0:0] comp_l1_p0_col12_cout;
	wire [0:0] comp_l1_p0_col12_sum ;
	wire [0:0] comp_l1_p0_col13_cout;
	wire [0:0] comp_l1_p0_col13_sum ;
	wire [0:0] comp_l1_p0_col14_cout;
	wire [0:0] comp_l1_p0_col14_sum ;
	wire [0:0] comp_l1_p0_col15_cout;
	wire [0:0] comp_l1_p0_col15_sum ;
	wire [0:0] comp_l1_p0_col16_cout;
	wire [0:0] comp_l1_p0_col16_sum ;
	wire [0:0] comp_l1_p0_col17_cout;
	wire [0:0] comp_l1_p0_col17_sum ;
	wire [0:0] comp_l1_p0_col18_cout;
	wire [0:0] comp_l1_p0_col18_sum ;
	wire [0:0] comp_l1_p0_col19_cout;
	wire [0:0] comp_l1_p0_col19_sum ;
	wire [0:0] comp_l1_p0_col20_cout;
	wire [0:0] comp_l1_p0_col20_sum ;
	wire [0:0] comp_l1_p0_col21_cout;
	wire [0:0] comp_l1_p0_col21_sum ;
	wire [0:0] comp_l1_p0_col22_cout;
	wire [0:0] comp_l1_p0_col22_sum ;
	wire [0:0] comp_l1_p0_col23_cout;
	wire [0:0] comp_l1_p0_col23_sum ;
	wire [0:0] comp_l1_p0_col24_cout;
	wire [0:0] comp_l1_p0_col24_sum ;
	wire [0:0] comp_l1_p0_col25_cout;
	wire [0:0] comp_l1_p0_col25_sum ;
	wire [0:0] comp_l1_p0_col26_cout;
	wire [0:0] comp_l1_p0_col26_sum ;
	wire [0:0] comp_l1_p0_col27_cout;
	wire [0:0] comp_l1_p0_col27_sum ;
	wire [0:0] comp_l1_p0_col28_cout;
	wire [0:0] comp_l1_p0_col28_sum ;
	wire [0:0] comp_l1_p0_col29_cout;
	wire [0:0] comp_l1_p0_col29_sum ;
	wire [0:0] comp_l1_p0_col30_cout;
	wire [0:0] comp_l1_p0_col30_sum ;
	wire [0:0] comp_l1_p0_col31_cout;
	wire [0:0] comp_l1_p0_col31_sum ;
	wire [0:0] comp_pad_l1_p0       ;
	wire [0:0] comp_l1_p1_col0_cout ;
	wire [0:0] comp_l1_p1_col0_sum  ;
	wire [0:0] comp_l1_p1_col1_cout ;
	wire [0:0] comp_l1_p1_col1_sum  ;
	wire [0:0] comp_l1_p1_col2_cout ;
	wire [0:0] comp_l1_p1_col2_sum  ;
	wire [0:0] comp_l1_p1_col3_cout ;
	wire [0:0] comp_l1_p1_col3_sum  ;
	wire [0:0] comp_l1_p1_col4_cout ;
	wire [0:0] comp_l1_p1_col4_sum  ;
	wire [0:0] comp_l1_p1_col5_cout ;
	wire [0:0] comp_l1_p1_col5_sum  ;
	wire [0:0] comp_l1_p1_col6_cout ;
	wire [0:0] comp_l1_p1_col6_sum  ;
	wire [0:0] comp_l1_p1_col7_cout ;
	wire [0:0] comp_l1_p1_col7_sum  ;
	wire [0:0] comp_l1_p1_col8_cout ;
	wire [0:0] comp_l1_p1_col8_sum  ;
	wire [0:0] comp_l1_p1_col9_cout ;
	wire [0:0] comp_l1_p1_col9_sum  ;
	wire [0:0] comp_l1_p1_col10_cout;
	wire [0:0] comp_l1_p1_col10_sum ;
	wire [0:0] comp_l1_p1_col11_cout;
	wire [0:0] comp_l1_p1_col11_sum ;
	wire [0:0] comp_l1_p1_col12_cout;
	wire [0:0] comp_l1_p1_col12_sum ;
	wire [0:0] comp_l1_p1_col13_cout;
	wire [0:0] comp_l1_p1_col13_sum ;
	wire [0:0] comp_l1_p1_col14_cout;
	wire [0:0] comp_l1_p1_col14_sum ;
	wire [0:0] comp_l1_p1_col15_cout;
	wire [0:0] comp_l1_p1_col15_sum ;
	wire [0:0] comp_l1_p1_col16_cout;
	wire [0:0] comp_l1_p1_col16_sum ;
	wire [0:0] comp_l1_p1_col17_cout;
	wire [0:0] comp_l1_p1_col17_sum ;
	wire [0:0] comp_l1_p1_col18_cout;
	wire [0:0] comp_l1_p1_col18_sum ;
	wire [0:0] comp_l1_p1_col19_cout;
	wire [0:0] comp_l1_p1_col19_sum ;
	wire [0:0] comp_l1_p1_col20_cout;
	wire [0:0] comp_l1_p1_col20_sum ;
	wire [0:0] comp_l1_p1_col21_cout;
	wire [0:0] comp_l1_p1_col21_sum ;
	wire [0:0] comp_l1_p1_col22_cout;
	wire [0:0] comp_l1_p1_col22_sum ;
	wire [0:0] comp_l1_p1_col23_cout;
	wire [0:0] comp_l1_p1_col23_sum ;
	wire [0:0] comp_l1_p1_col24_cout;
	wire [0:0] comp_l1_p1_col24_sum ;
	wire [0:0] comp_l1_p1_col25_cout;
	wire [0:0] comp_l1_p1_col25_sum ;
	wire [0:0] comp_l1_p1_col26_cout;
	wire [0:0] comp_l1_p1_col26_sum ;
	wire [0:0] comp_l1_p1_col27_cout;
	wire [0:0] comp_l1_p1_col27_sum ;
	wire [0:0] comp_l1_p1_col28_cout;
	wire [0:0] comp_l1_p1_col28_sum ;
	wire [0:0] comp_l1_p1_col29_cout;
	wire [0:0] comp_l1_p1_col29_sum ;
	wire [0:0] comp_l1_p1_col30_cout;
	wire [0:0] comp_l1_p1_col30_sum ;
	wire [0:0] comp_l1_p1_col31_cout;
	wire [0:0] comp_l1_p1_col31_sum ;
	wire [0:0] comp_pad_l1_p1       ;
	wire [0:0] comp_l2_p0_col0_cout ;
	wire [0:0] comp_l2_p0_col0_sum  ;
	wire [0:0] comp_l2_p0_col1_cout ;
	wire [0:0] comp_l2_p0_col1_sum  ;
	wire [0:0] comp_l2_p0_col2_cout ;
	wire [0:0] comp_l2_p0_col2_sum  ;
	wire [0:0] comp_l2_p0_col3_cout ;
	wire [0:0] comp_l2_p0_col3_sum  ;
	wire [0:0] comp_l2_p0_col4_cout ;
	wire [0:0] comp_l2_p0_col4_sum  ;
	wire [0:0] comp_l2_p0_col5_cout ;
	wire [0:0] comp_l2_p0_col5_sum  ;
	wire [0:0] comp_l2_p0_col6_cout ;
	wire [0:0] comp_l2_p0_col6_sum  ;
	wire [0:0] comp_l2_p0_col7_cout ;
	wire [0:0] comp_l2_p0_col7_sum  ;
	wire [0:0] comp_l2_p0_col8_cout ;
	wire [0:0] comp_l2_p0_col8_sum  ;
	wire [0:0] comp_l2_p0_col9_cout ;
	wire [0:0] comp_l2_p0_col9_sum  ;
	wire [0:0] comp_l2_p0_col10_cout;
	wire [0:0] comp_l2_p0_col10_sum ;
	wire [0:0] comp_l2_p0_col11_cout;
	wire [0:0] comp_l2_p0_col11_sum ;
	wire [0:0] comp_l2_p0_col12_cout;
	wire [0:0] comp_l2_p0_col12_sum ;
	wire [0:0] comp_l2_p0_col13_cout;
	wire [0:0] comp_l2_p0_col13_sum ;
	wire [0:0] comp_l2_p0_col14_cout;
	wire [0:0] comp_l2_p0_col14_sum ;
	wire [0:0] comp_l2_p0_col15_cout;
	wire [0:0] comp_l2_p0_col15_sum ;
	wire [0:0] comp_l2_p0_col16_cout;
	wire [0:0] comp_l2_p0_col16_sum ;
	wire [0:0] comp_l2_p0_col17_cout;
	wire [0:0] comp_l2_p0_col17_sum ;
	wire [0:0] comp_l2_p0_col18_cout;
	wire [0:0] comp_l2_p0_col18_sum ;
	wire [0:0] comp_l2_p0_col19_cout;
	wire [0:0] comp_l2_p0_col19_sum ;
	wire [0:0] comp_l2_p0_col20_cout;
	wire [0:0] comp_l2_p0_col20_sum ;
	wire [0:0] comp_l2_p0_col21_cout;
	wire [0:0] comp_l2_p0_col21_sum ;
	wire [0:0] comp_l2_p0_col22_cout;
	wire [0:0] comp_l2_p0_col22_sum ;
	wire [0:0] comp_l2_p0_col23_cout;
	wire [0:0] comp_l2_p0_col23_sum ;
	wire [0:0] comp_l2_p0_col24_cout;
	wire [0:0] comp_l2_p0_col24_sum ;
	wire [0:0] comp_l2_p0_col25_cout;
	wire [0:0] comp_l2_p0_col25_sum ;
	wire [0:0] comp_l2_p0_col26_cout;
	wire [0:0] comp_l2_p0_col26_sum ;
	wire [0:0] comp_l2_p0_col27_cout;
	wire [0:0] comp_l2_p0_col27_sum ;
	wire [0:0] comp_l2_p0_col28_cout;
	wire [0:0] comp_l2_p0_col28_sum ;
	wire [0:0] comp_l2_p0_col29_cout;
	wire [0:0] comp_l2_p0_col29_sum ;
	wire [0:0] comp_l2_p0_col30_cout;
	wire [0:0] comp_l2_p0_col30_sum ;
	wire [0:0] comp_l2_p0_col31_cout;
	wire [0:0] comp_l2_p0_col31_sum ;
	wire [0:0] comp_pad_l2_p0       ;
	wire [0:0] comp_l3_p0_col0_cout ;
	wire [0:0] comp_l3_p0_col0_sum  ;
	wire [0:0] comp_l3_p0_col1_cout ;
	wire [0:0] comp_l3_p0_col1_sum  ;
	wire [0:0] comp_l3_p0_col2_cout ;
	wire [0:0] comp_l3_p0_col2_sum  ;
	wire [0:0] comp_l3_p0_col3_cout ;
	wire [0:0] comp_l3_p0_col3_sum  ;
	wire [0:0] comp_l3_p0_col4_cout ;
	wire [0:0] comp_l3_p0_col4_sum  ;
	wire [0:0] comp_l3_p0_col5_cout ;
	wire [0:0] comp_l3_p0_col5_sum  ;
	wire [0:0] comp_l3_p0_col6_cout ;
	wire [0:0] comp_l3_p0_col6_sum  ;
	wire [0:0] comp_l3_p0_col7_cout ;
	wire [0:0] comp_l3_p0_col7_sum  ;
	wire [0:0] comp_l3_p0_col8_cout ;
	wire [0:0] comp_l3_p0_col8_sum  ;
	wire [0:0] comp_l3_p0_col9_cout ;
	wire [0:0] comp_l3_p0_col9_sum  ;
	wire [0:0] comp_l3_p0_col10_cout;
	wire [0:0] comp_l3_p0_col10_sum ;
	wire [0:0] comp_l3_p0_col11_cout;
	wire [0:0] comp_l3_p0_col11_sum ;
	wire [0:0] comp_l3_p0_col12_cout;
	wire [0:0] comp_l3_p0_col12_sum ;
	wire [0:0] comp_l3_p0_col13_cout;
	wire [0:0] comp_l3_p0_col13_sum ;
	wire [0:0] comp_l3_p0_col14_cout;
	wire [0:0] comp_l3_p0_col14_sum ;
	wire [0:0] comp_l3_p0_col15_cout;
	wire [0:0] comp_l3_p0_col15_sum ;
	wire [0:0] comp_l3_p0_col16_cout;
	wire [0:0] comp_l3_p0_col16_sum ;
	wire [0:0] comp_l3_p0_col17_cout;
	wire [0:0] comp_l3_p0_col17_sum ;
	wire [0:0] comp_l3_p0_col18_cout;
	wire [0:0] comp_l3_p0_col18_sum ;
	wire [0:0] comp_l3_p0_col19_cout;
	wire [0:0] comp_l3_p0_col19_sum ;
	wire [0:0] comp_l3_p0_col20_cout;
	wire [0:0] comp_l3_p0_col20_sum ;
	wire [0:0] comp_l3_p0_col21_cout;
	wire [0:0] comp_l3_p0_col21_sum ;
	wire [0:0] comp_l3_p0_col22_cout;
	wire [0:0] comp_l3_p0_col22_sum ;
	wire [0:0] comp_l3_p0_col23_cout;
	wire [0:0] comp_l3_p0_col23_sum ;
	wire [0:0] comp_l3_p0_col24_cout;
	wire [0:0] comp_l3_p0_col24_sum ;
	wire [0:0] comp_l3_p0_col25_cout;
	wire [0:0] comp_l3_p0_col25_sum ;
	wire [0:0] comp_l3_p0_col26_cout;
	wire [0:0] comp_l3_p0_col26_sum ;
	wire [0:0] comp_l3_p0_col27_cout;
	wire [0:0] comp_l3_p0_col27_sum ;
	wire [0:0] comp_l3_p0_col28_cout;
	wire [0:0] comp_l3_p0_col28_sum ;
	wire [0:0] comp_l3_p0_col29_cout;
	wire [0:0] comp_l3_p0_col29_sum ;
	wire [0:0] comp_l3_p0_col30_cout;
	wire [0:0] comp_l3_p0_col30_sum ;
	wire [0:0] comp_l3_p0_col31_cout;
	wire [0:0] comp_l3_p0_col31_sum ;
	wire [0:0] comp_pad_l3_p0       ;
	wire [0:0] comp_l4_p0_col0_cout ;
	wire [0:0] comp_l4_p0_col0_sum  ;
	wire [0:0] comp_l4_p0_col1_cout ;
	wire [0:0] comp_l4_p0_col1_sum  ;
	wire [0:0] comp_l4_p0_col2_cout ;
	wire [0:0] comp_l4_p0_col2_sum  ;
	wire [0:0] comp_l4_p0_col3_cout ;
	wire [0:0] comp_l4_p0_col3_sum  ;
	wire [0:0] comp_l4_p0_col4_cout ;
	wire [0:0] comp_l4_p0_col4_sum  ;
	wire [0:0] comp_l4_p0_col5_cout ;
	wire [0:0] comp_l4_p0_col5_sum  ;
	wire [0:0] comp_l4_p0_col6_cout ;
	wire [0:0] comp_l4_p0_col6_sum  ;
	wire [0:0] comp_l4_p0_col7_cout ;
	wire [0:0] comp_l4_p0_col7_sum  ;
	wire [0:0] comp_l4_p0_col8_cout ;
	wire [0:0] comp_l4_p0_col8_sum  ;
	wire [0:0] comp_l4_p0_col9_cout ;
	wire [0:0] comp_l4_p0_col9_sum  ;
	wire [0:0] comp_l4_p0_col10_cout;
	wire [0:0] comp_l4_p0_col10_sum ;
	wire [0:0] comp_l4_p0_col11_cout;
	wire [0:0] comp_l4_p0_col11_sum ;
	wire [0:0] comp_l4_p0_col12_cout;
	wire [0:0] comp_l4_p0_col12_sum ;
	wire [0:0] comp_l4_p0_col13_cout;
	wire [0:0] comp_l4_p0_col13_sum ;
	wire [0:0] comp_l4_p0_col14_cout;
	wire [0:0] comp_l4_p0_col14_sum ;
	wire [0:0] comp_l4_p0_col15_cout;
	wire [0:0] comp_l4_p0_col15_sum ;
	wire [0:0] comp_l4_p0_col16_cout;
	wire [0:0] comp_l4_p0_col16_sum ;
	wire [0:0] comp_l4_p0_col17_cout;
	wire [0:0] comp_l4_p0_col17_sum ;
	wire [0:0] comp_l4_p0_col18_cout;
	wire [0:0] comp_l4_p0_col18_sum ;
	wire [0:0] comp_l4_p0_col19_cout;
	wire [0:0] comp_l4_p0_col19_sum ;
	wire [0:0] comp_l4_p0_col20_cout;
	wire [0:0] comp_l4_p0_col20_sum ;
	wire [0:0] comp_l4_p0_col21_cout;
	wire [0:0] comp_l4_p0_col21_sum ;
	wire [0:0] comp_l4_p0_col22_cout;
	wire [0:0] comp_l4_p0_col22_sum ;
	wire [0:0] comp_l4_p0_col23_cout;
	wire [0:0] comp_l4_p0_col23_sum ;
	wire [0:0] comp_l4_p0_col24_cout;
	wire [0:0] comp_l4_p0_col24_sum ;
	wire [0:0] comp_l4_p0_col25_cout;
	wire [0:0] comp_l4_p0_col25_sum ;
	wire [0:0] comp_l4_p0_col26_cout;
	wire [0:0] comp_l4_p0_col26_sum ;
	wire [0:0] comp_l4_p0_col27_cout;
	wire [0:0] comp_l4_p0_col27_sum ;
	wire [0:0] comp_l4_p0_col28_cout;
	wire [0:0] comp_l4_p0_col28_sum ;
	wire [0:0] comp_l4_p0_col29_cout;
	wire [0:0] comp_l4_p0_col29_sum ;
	wire [0:0] comp_l4_p0_col30_cout;
	wire [0:0] comp_l4_p0_col30_sum ;
	wire [0:0] comp_l4_p0_col31_cout;
	wire [0:0] comp_l4_p0_col31_sum ;
	wire [0:0] comp_pad_l4_p0       ;

	//Wire define for sub module.
	wire  u_comp_l0_p0_col0_cout ;
	wire  u_comp_l0_p0_col0_sum  ;
	wire  u_comp_l0_p0_col1_cout ;
	wire  u_comp_l0_p0_col1_sum  ;
	wire  u_comp_l0_p0_col2_cout ;
	wire  u_comp_l0_p0_col2_sum  ;
	wire  u_comp_l0_p0_col3_cout ;
	wire  u_comp_l0_p0_col3_sum  ;
	wire  u_comp_l0_p0_col4_cout ;
	wire  u_comp_l0_p0_col4_sum  ;
	wire  u_comp_l0_p0_col5_cout ;
	wire  u_comp_l0_p0_col5_sum  ;
	wire  u_comp_l0_p0_col6_cout ;
	wire  u_comp_l0_p0_col6_sum  ;
	wire  u_comp_l0_p0_col7_cout ;
	wire  u_comp_l0_p0_col7_sum  ;
	wire  u_comp_l0_p0_col8_cout ;
	wire  u_comp_l0_p0_col8_sum  ;
	wire  u_comp_l0_p0_col9_cout ;
	wire  u_comp_l0_p0_col9_sum  ;
	wire  u_comp_l0_p0_col10_cout;
	wire  u_comp_l0_p0_col10_sum ;
	wire  u_comp_l0_p0_col11_cout;
	wire  u_comp_l0_p0_col11_sum ;
	wire  u_comp_l0_p0_col12_cout;
	wire  u_comp_l0_p0_col12_sum ;
	wire  u_comp_l0_p0_col13_cout;
	wire  u_comp_l0_p0_col13_sum ;
	wire  u_comp_l0_p0_col14_cout;
	wire  u_comp_l0_p0_col14_sum ;
	wire  u_comp_l0_p0_col15_cout;
	wire  u_comp_l0_p0_col15_sum ;
	wire  u_comp_l0_p0_col16_cout;
	wire  u_comp_l0_p0_col16_sum ;
	wire  u_comp_l0_p0_col17_cout;
	wire  u_comp_l0_p0_col17_sum ;
	wire  u_comp_l0_p0_col18_cout;
	wire  u_comp_l0_p0_col18_sum ;
	wire  u_comp_l0_p0_col19_cout;
	wire  u_comp_l0_p0_col19_sum ;
	wire  u_comp_l0_p0_col20_cout;
	wire  u_comp_l0_p0_col20_sum ;
	wire  u_comp_l0_p0_col21_cout;
	wire  u_comp_l0_p0_col21_sum ;
	wire  u_comp_l0_p0_col22_cout;
	wire  u_comp_l0_p0_col22_sum ;
	wire  u_comp_l0_p0_col23_cout;
	wire  u_comp_l0_p0_col23_sum ;
	wire  u_comp_l0_p0_col24_cout;
	wire  u_comp_l0_p0_col24_sum ;
	wire  u_comp_l0_p0_col25_cout;
	wire  u_comp_l0_p0_col25_sum ;
	wire  u_comp_l0_p0_col26_cout;
	wire  u_comp_l0_p0_col26_sum ;
	wire  u_comp_l0_p0_col27_cout;
	wire  u_comp_l0_p0_col27_sum ;
	wire  u_comp_l0_p0_col28_cout;
	wire  u_comp_l0_p0_col28_sum ;
	wire  u_comp_l0_p0_col29_cout;
	wire  u_comp_l0_p0_col29_sum ;
	wire  u_comp_l0_p0_col30_cout;
	wire  u_comp_l0_p0_col30_sum ;
	wire  u_comp_l0_p0_col31_sum ;
	wire  u_comp_l0_p1_col0_cout ;
	wire  u_comp_l0_p1_col0_sum  ;
	wire  u_comp_l0_p1_col1_cout ;
	wire  u_comp_l0_p1_col1_sum  ;
	wire  u_comp_l0_p1_col2_cout ;
	wire  u_comp_l0_p1_col2_sum  ;
	wire  u_comp_l0_p1_col3_cout ;
	wire  u_comp_l0_p1_col3_sum  ;
	wire  u_comp_l0_p1_col4_cout ;
	wire  u_comp_l0_p1_col4_sum  ;
	wire  u_comp_l0_p1_col5_cout ;
	wire  u_comp_l0_p1_col5_sum  ;
	wire  u_comp_l0_p1_col6_cout ;
	wire  u_comp_l0_p1_col6_sum  ;
	wire  u_comp_l0_p1_col7_cout ;
	wire  u_comp_l0_p1_col7_sum  ;
	wire  u_comp_l0_p1_col8_cout ;
	wire  u_comp_l0_p1_col8_sum  ;
	wire  u_comp_l0_p1_col9_cout ;
	wire  u_comp_l0_p1_col9_sum  ;
	wire  u_comp_l0_p1_col10_cout;
	wire  u_comp_l0_p1_col10_sum ;
	wire  u_comp_l0_p1_col11_cout;
	wire  u_comp_l0_p1_col11_sum ;
	wire  u_comp_l0_p1_col12_cout;
	wire  u_comp_l0_p1_col12_sum ;
	wire  u_comp_l0_p1_col13_cout;
	wire  u_comp_l0_p1_col13_sum ;
	wire  u_comp_l0_p1_col14_cout;
	wire  u_comp_l0_p1_col14_sum ;
	wire  u_comp_l0_p1_col15_cout;
	wire  u_comp_l0_p1_col15_sum ;
	wire  u_comp_l0_p1_col16_cout;
	wire  u_comp_l0_p1_col16_sum ;
	wire  u_comp_l0_p1_col17_cout;
	wire  u_comp_l0_p1_col17_sum ;
	wire  u_comp_l0_p1_col18_cout;
	wire  u_comp_l0_p1_col18_sum ;
	wire  u_comp_l0_p1_col19_cout;
	wire  u_comp_l0_p1_col19_sum ;
	wire  u_comp_l0_p1_col20_cout;
	wire  u_comp_l0_p1_col20_sum ;
	wire  u_comp_l0_p1_col21_cout;
	wire  u_comp_l0_p1_col21_sum ;
	wire  u_comp_l0_p1_col22_cout;
	wire  u_comp_l0_p1_col22_sum ;
	wire  u_comp_l0_p1_col23_cout;
	wire  u_comp_l0_p1_col23_sum ;
	wire  u_comp_l0_p1_col24_cout;
	wire  u_comp_l0_p1_col24_sum ;
	wire  u_comp_l0_p1_col25_cout;
	wire  u_comp_l0_p1_col25_sum ;
	wire  u_comp_l0_p1_col26_cout;
	wire  u_comp_l0_p1_col26_sum ;
	wire  u_comp_l0_p1_col27_cout;
	wire  u_comp_l0_p1_col27_sum ;
	wire  u_comp_l0_p1_col28_cout;
	wire  u_comp_l0_p1_col28_sum ;
	wire  u_comp_l0_p1_col29_cout;
	wire  u_comp_l0_p1_col29_sum ;
	wire  u_comp_l0_p1_col30_cout;
	wire  u_comp_l0_p1_col30_sum ;
	wire  u_comp_l0_p1_col31_sum ;
	wire  u_comp_l0_p2_col0_cout ;
	wire  u_comp_l0_p2_col0_sum  ;
	wire  u_comp_l0_p2_col1_cout ;
	wire  u_comp_l0_p2_col1_sum  ;
	wire  u_comp_l0_p2_col2_cout ;
	wire  u_comp_l0_p2_col2_sum  ;
	wire  u_comp_l0_p2_col3_cout ;
	wire  u_comp_l0_p2_col3_sum  ;
	wire  u_comp_l0_p2_col4_cout ;
	wire  u_comp_l0_p2_col4_sum  ;
	wire  u_comp_l0_p2_col5_cout ;
	wire  u_comp_l0_p2_col5_sum  ;
	wire  u_comp_l0_p2_col6_cout ;
	wire  u_comp_l0_p2_col6_sum  ;
	wire  u_comp_l0_p2_col7_cout ;
	wire  u_comp_l0_p2_col7_sum  ;
	wire  u_comp_l0_p2_col8_cout ;
	wire  u_comp_l0_p2_col8_sum  ;
	wire  u_comp_l0_p2_col9_cout ;
	wire  u_comp_l0_p2_col9_sum  ;
	wire  u_comp_l0_p2_col10_cout;
	wire  u_comp_l0_p2_col10_sum ;
	wire  u_comp_l0_p2_col11_cout;
	wire  u_comp_l0_p2_col11_sum ;
	wire  u_comp_l0_p2_col12_cout;
	wire  u_comp_l0_p2_col12_sum ;
	wire  u_comp_l0_p2_col13_cout;
	wire  u_comp_l0_p2_col13_sum ;
	wire  u_comp_l0_p2_col14_cout;
	wire  u_comp_l0_p2_col14_sum ;
	wire  u_comp_l0_p2_col15_cout;
	wire  u_comp_l0_p2_col15_sum ;
	wire  u_comp_l0_p2_col16_cout;
	wire  u_comp_l0_p2_col16_sum ;
	wire  u_comp_l0_p2_col17_cout;
	wire  u_comp_l0_p2_col17_sum ;
	wire  u_comp_l0_p2_col18_cout;
	wire  u_comp_l0_p2_col18_sum ;
	wire  u_comp_l0_p2_col19_cout;
	wire  u_comp_l0_p2_col19_sum ;
	wire  u_comp_l0_p2_col20_cout;
	wire  u_comp_l0_p2_col20_sum ;
	wire  u_comp_l0_p2_col21_cout;
	wire  u_comp_l0_p2_col21_sum ;
	wire  u_comp_l0_p2_col22_cout;
	wire  u_comp_l0_p2_col22_sum ;
	wire  u_comp_l0_p2_col23_cout;
	wire  u_comp_l0_p2_col23_sum ;
	wire  u_comp_l0_p2_col24_cout;
	wire  u_comp_l0_p2_col24_sum ;
	wire  u_comp_l0_p2_col25_cout;
	wire  u_comp_l0_p2_col25_sum ;
	wire  u_comp_l0_p2_col26_cout;
	wire  u_comp_l0_p2_col26_sum ;
	wire  u_comp_l0_p2_col27_cout;
	wire  u_comp_l0_p2_col27_sum ;
	wire  u_comp_l0_p2_col28_cout;
	wire  u_comp_l0_p2_col28_sum ;
	wire  u_comp_l0_p2_col29_cout;
	wire  u_comp_l0_p2_col29_sum ;
	wire  u_comp_l0_p2_col30_cout;
	wire  u_comp_l0_p2_col30_sum ;
	wire  u_comp_l0_p2_col31_sum ;
	wire  u_comp_l1_p0_col0_cout ;
	wire  u_comp_l1_p0_col0_sum  ;
	wire  u_comp_l1_p0_col1_cout ;
	wire  u_comp_l1_p0_col1_sum  ;
	wire  u_comp_l1_p0_col2_cout ;
	wire  u_comp_l1_p0_col2_sum  ;
	wire  u_comp_l1_p0_col3_cout ;
	wire  u_comp_l1_p0_col3_sum  ;
	wire  u_comp_l1_p0_col4_cout ;
	wire  u_comp_l1_p0_col4_sum  ;
	wire  u_comp_l1_p0_col5_cout ;
	wire  u_comp_l1_p0_col5_sum  ;
	wire  u_comp_l1_p0_col6_cout ;
	wire  u_comp_l1_p0_col6_sum  ;
	wire  u_comp_l1_p0_col7_cout ;
	wire  u_comp_l1_p0_col7_sum  ;
	wire  u_comp_l1_p0_col8_cout ;
	wire  u_comp_l1_p0_col8_sum  ;
	wire  u_comp_l1_p0_col9_cout ;
	wire  u_comp_l1_p0_col9_sum  ;
	wire  u_comp_l1_p0_col10_cout;
	wire  u_comp_l1_p0_col10_sum ;
	wire  u_comp_l1_p0_col11_cout;
	wire  u_comp_l1_p0_col11_sum ;
	wire  u_comp_l1_p0_col12_cout;
	wire  u_comp_l1_p0_col12_sum ;
	wire  u_comp_l1_p0_col13_cout;
	wire  u_comp_l1_p0_col13_sum ;
	wire  u_comp_l1_p0_col14_cout;
	wire  u_comp_l1_p0_col14_sum ;
	wire  u_comp_l1_p0_col15_cout;
	wire  u_comp_l1_p0_col15_sum ;
	wire  u_comp_l1_p0_col16_cout;
	wire  u_comp_l1_p0_col16_sum ;
	wire  u_comp_l1_p0_col17_cout;
	wire  u_comp_l1_p0_col17_sum ;
	wire  u_comp_l1_p0_col18_cout;
	wire  u_comp_l1_p0_col18_sum ;
	wire  u_comp_l1_p0_col19_cout;
	wire  u_comp_l1_p0_col19_sum ;
	wire  u_comp_l1_p0_col20_cout;
	wire  u_comp_l1_p0_col20_sum ;
	wire  u_comp_l1_p0_col21_cout;
	wire  u_comp_l1_p0_col21_sum ;
	wire  u_comp_l1_p0_col22_cout;
	wire  u_comp_l1_p0_col22_sum ;
	wire  u_comp_l1_p0_col23_cout;
	wire  u_comp_l1_p0_col23_sum ;
	wire  u_comp_l1_p0_col24_cout;
	wire  u_comp_l1_p0_col24_sum ;
	wire  u_comp_l1_p0_col25_cout;
	wire  u_comp_l1_p0_col25_sum ;
	wire  u_comp_l1_p0_col26_cout;
	wire  u_comp_l1_p0_col26_sum ;
	wire  u_comp_l1_p0_col27_cout;
	wire  u_comp_l1_p0_col27_sum ;
	wire  u_comp_l1_p0_col28_cout;
	wire  u_comp_l1_p0_col28_sum ;
	wire  u_comp_l1_p0_col29_cout;
	wire  u_comp_l1_p0_col29_sum ;
	wire  u_comp_l1_p0_col30_cout;
	wire  u_comp_l1_p0_col30_sum ;
	wire  u_comp_l1_p0_col31_sum ;
	wire  u_comp_l1_p1_col0_cout ;
	wire  u_comp_l1_p1_col0_sum  ;
	wire  u_comp_l1_p1_col1_cout ;
	wire  u_comp_l1_p1_col1_sum  ;
	wire  u_comp_l1_p1_col2_cout ;
	wire  u_comp_l1_p1_col2_sum  ;
	wire  u_comp_l1_p1_col3_cout ;
	wire  u_comp_l1_p1_col3_sum  ;
	wire  u_comp_l1_p1_col4_cout ;
	wire  u_comp_l1_p1_col4_sum  ;
	wire  u_comp_l1_p1_col5_cout ;
	wire  u_comp_l1_p1_col5_sum  ;
	wire  u_comp_l1_p1_col6_cout ;
	wire  u_comp_l1_p1_col6_sum  ;
	wire  u_comp_l1_p1_col7_cout ;
	wire  u_comp_l1_p1_col7_sum  ;
	wire  u_comp_l1_p1_col8_cout ;
	wire  u_comp_l1_p1_col8_sum  ;
	wire  u_comp_l1_p1_col9_cout ;
	wire  u_comp_l1_p1_col9_sum  ;
	wire  u_comp_l1_p1_col10_cout;
	wire  u_comp_l1_p1_col10_sum ;
	wire  u_comp_l1_p1_col11_cout;
	wire  u_comp_l1_p1_col11_sum ;
	wire  u_comp_l1_p1_col12_cout;
	wire  u_comp_l1_p1_col12_sum ;
	wire  u_comp_l1_p1_col13_cout;
	wire  u_comp_l1_p1_col13_sum ;
	wire  u_comp_l1_p1_col14_cout;
	wire  u_comp_l1_p1_col14_sum ;
	wire  u_comp_l1_p1_col15_cout;
	wire  u_comp_l1_p1_col15_sum ;
	wire  u_comp_l1_p1_col16_cout;
	wire  u_comp_l1_p1_col16_sum ;
	wire  u_comp_l1_p1_col17_cout;
	wire  u_comp_l1_p1_col17_sum ;
	wire  u_comp_l1_p1_col18_cout;
	wire  u_comp_l1_p1_col18_sum ;
	wire  u_comp_l1_p1_col19_cout;
	wire  u_comp_l1_p1_col19_sum ;
	wire  u_comp_l1_p1_col20_cout;
	wire  u_comp_l1_p1_col20_sum ;
	wire  u_comp_l1_p1_col21_cout;
	wire  u_comp_l1_p1_col21_sum ;
	wire  u_comp_l1_p1_col22_cout;
	wire  u_comp_l1_p1_col22_sum ;
	wire  u_comp_l1_p1_col23_cout;
	wire  u_comp_l1_p1_col23_sum ;
	wire  u_comp_l1_p1_col24_cout;
	wire  u_comp_l1_p1_col24_sum ;
	wire  u_comp_l1_p1_col25_cout;
	wire  u_comp_l1_p1_col25_sum ;
	wire  u_comp_l1_p1_col26_cout;
	wire  u_comp_l1_p1_col26_sum ;
	wire  u_comp_l1_p1_col27_cout;
	wire  u_comp_l1_p1_col27_sum ;
	wire  u_comp_l1_p1_col28_cout;
	wire  u_comp_l1_p1_col28_sum ;
	wire  u_comp_l1_p1_col29_cout;
	wire  u_comp_l1_p1_col29_sum ;
	wire  u_comp_l1_p1_col30_cout;
	wire  u_comp_l1_p1_col30_sum ;
	wire  u_comp_l1_p1_col31_sum ;
	wire  u_comp_l2_p0_col0_cout ;
	wire  u_comp_l2_p0_col0_sum  ;
	wire  u_comp_l2_p0_col1_cout ;
	wire  u_comp_l2_p0_col1_sum  ;
	wire  u_comp_l2_p0_col2_cout ;
	wire  u_comp_l2_p0_col2_sum  ;
	wire  u_comp_l2_p0_col3_cout ;
	wire  u_comp_l2_p0_col3_sum  ;
	wire  u_comp_l2_p0_col4_cout ;
	wire  u_comp_l2_p0_col4_sum  ;
	wire  u_comp_l2_p0_col5_cout ;
	wire  u_comp_l2_p0_col5_sum  ;
	wire  u_comp_l2_p0_col6_cout ;
	wire  u_comp_l2_p0_col6_sum  ;
	wire  u_comp_l2_p0_col7_cout ;
	wire  u_comp_l2_p0_col7_sum  ;
	wire  u_comp_l2_p0_col8_cout ;
	wire  u_comp_l2_p0_col8_sum  ;
	wire  u_comp_l2_p0_col9_cout ;
	wire  u_comp_l2_p0_col9_sum  ;
	wire  u_comp_l2_p0_col10_cout;
	wire  u_comp_l2_p0_col10_sum ;
	wire  u_comp_l2_p0_col11_cout;
	wire  u_comp_l2_p0_col11_sum ;
	wire  u_comp_l2_p0_col12_cout;
	wire  u_comp_l2_p0_col12_sum ;
	wire  u_comp_l2_p0_col13_cout;
	wire  u_comp_l2_p0_col13_sum ;
	wire  u_comp_l2_p0_col14_cout;
	wire  u_comp_l2_p0_col14_sum ;
	wire  u_comp_l2_p0_col15_cout;
	wire  u_comp_l2_p0_col15_sum ;
	wire  u_comp_l2_p0_col16_cout;
	wire  u_comp_l2_p0_col16_sum ;
	wire  u_comp_l2_p0_col17_cout;
	wire  u_comp_l2_p0_col17_sum ;
	wire  u_comp_l2_p0_col18_cout;
	wire  u_comp_l2_p0_col18_sum ;
	wire  u_comp_l2_p0_col19_cout;
	wire  u_comp_l2_p0_col19_sum ;
	wire  u_comp_l2_p0_col20_cout;
	wire  u_comp_l2_p0_col20_sum ;
	wire  u_comp_l2_p0_col21_cout;
	wire  u_comp_l2_p0_col21_sum ;
	wire  u_comp_l2_p0_col22_cout;
	wire  u_comp_l2_p0_col22_sum ;
	wire  u_comp_l2_p0_col23_cout;
	wire  u_comp_l2_p0_col23_sum ;
	wire  u_comp_l2_p0_col24_cout;
	wire  u_comp_l2_p0_col24_sum ;
	wire  u_comp_l2_p0_col25_cout;
	wire  u_comp_l2_p0_col25_sum ;
	wire  u_comp_l2_p0_col26_cout;
	wire  u_comp_l2_p0_col26_sum ;
	wire  u_comp_l2_p0_col27_cout;
	wire  u_comp_l2_p0_col27_sum ;
	wire  u_comp_l2_p0_col28_cout;
	wire  u_comp_l2_p0_col28_sum ;
	wire  u_comp_l2_p0_col29_cout;
	wire  u_comp_l2_p0_col29_sum ;
	wire  u_comp_l2_p0_col30_cout;
	wire  u_comp_l2_p0_col30_sum ;
	wire  u_comp_l2_p0_col31_sum ;
	wire  u_comp_l3_p0_col0_cout ;
	wire  u_comp_l3_p0_col0_sum  ;
	wire  u_comp_l3_p0_col1_cout ;
	wire  u_comp_l3_p0_col1_sum  ;
	wire  u_comp_l3_p0_col2_cout ;
	wire  u_comp_l3_p0_col2_sum  ;
	wire  u_comp_l3_p0_col3_cout ;
	wire  u_comp_l3_p0_col3_sum  ;
	wire  u_comp_l3_p0_col4_cout ;
	wire  u_comp_l3_p0_col4_sum  ;
	wire  u_comp_l3_p0_col5_cout ;
	wire  u_comp_l3_p0_col5_sum  ;
	wire  u_comp_l3_p0_col6_cout ;
	wire  u_comp_l3_p0_col6_sum  ;
	wire  u_comp_l3_p0_col7_cout ;
	wire  u_comp_l3_p0_col7_sum  ;
	wire  u_comp_l3_p0_col8_cout ;
	wire  u_comp_l3_p0_col8_sum  ;
	wire  u_comp_l3_p0_col9_cout ;
	wire  u_comp_l3_p0_col9_sum  ;
	wire  u_comp_l3_p0_col10_cout;
	wire  u_comp_l3_p0_col10_sum ;
	wire  u_comp_l3_p0_col11_cout;
	wire  u_comp_l3_p0_col11_sum ;
	wire  u_comp_l3_p0_col12_cout;
	wire  u_comp_l3_p0_col12_sum ;
	wire  u_comp_l3_p0_col13_cout;
	wire  u_comp_l3_p0_col13_sum ;
	wire  u_comp_l3_p0_col14_cout;
	wire  u_comp_l3_p0_col14_sum ;
	wire  u_comp_l3_p0_col15_cout;
	wire  u_comp_l3_p0_col15_sum ;
	wire  u_comp_l3_p0_col16_cout;
	wire  u_comp_l3_p0_col16_sum ;
	wire  u_comp_l3_p0_col17_cout;
	wire  u_comp_l3_p0_col17_sum ;
	wire  u_comp_l3_p0_col18_cout;
	wire  u_comp_l3_p0_col18_sum ;
	wire  u_comp_l3_p0_col19_cout;
	wire  u_comp_l3_p0_col19_sum ;
	wire  u_comp_l3_p0_col20_cout;
	wire  u_comp_l3_p0_col20_sum ;
	wire  u_comp_l3_p0_col21_cout;
	wire  u_comp_l3_p0_col21_sum ;
	wire  u_comp_l3_p0_col22_cout;
	wire  u_comp_l3_p0_col22_sum ;
	wire  u_comp_l3_p0_col23_cout;
	wire  u_comp_l3_p0_col23_sum ;
	wire  u_comp_l3_p0_col24_cout;
	wire  u_comp_l3_p0_col24_sum ;
	wire  u_comp_l3_p0_col25_cout;
	wire  u_comp_l3_p0_col25_sum ;
	wire  u_comp_l3_p0_col26_cout;
	wire  u_comp_l3_p0_col26_sum ;
	wire  u_comp_l3_p0_col27_cout;
	wire  u_comp_l3_p0_col27_sum ;
	wire  u_comp_l3_p0_col28_cout;
	wire  u_comp_l3_p0_col28_sum ;
	wire  u_comp_l3_p0_col29_cout;
	wire  u_comp_l3_p0_col29_sum ;
	wire  u_comp_l3_p0_col30_cout;
	wire  u_comp_l3_p0_col30_sum ;
	wire  u_comp_l3_p0_col31_sum ;
	wire  u_comp_l4_p0_col0_cout ;
	wire  u_comp_l4_p0_col0_sum  ;
	wire  u_comp_l4_p0_col1_cout ;
	wire  u_comp_l4_p0_col1_sum  ;
	wire  u_comp_l4_p0_col2_cout ;
	wire  u_comp_l4_p0_col2_sum  ;
	wire  u_comp_l4_p0_col3_cout ;
	wire  u_comp_l4_p0_col3_sum  ;
	wire  u_comp_l4_p0_col4_cout ;
	wire  u_comp_l4_p0_col4_sum  ;
	wire  u_comp_l4_p0_col5_cout ;
	wire  u_comp_l4_p0_col5_sum  ;
	wire  u_comp_l4_p0_col6_cout ;
	wire  u_comp_l4_p0_col6_sum  ;
	wire  u_comp_l4_p0_col7_cout ;
	wire  u_comp_l4_p0_col7_sum  ;
	wire  u_comp_l4_p0_col8_cout ;
	wire  u_comp_l4_p0_col8_sum  ;
	wire  u_comp_l4_p0_col9_cout ;
	wire  u_comp_l4_p0_col9_sum  ;
	wire  u_comp_l4_p0_col10_cout;
	wire  u_comp_l4_p0_col10_sum ;
	wire  u_comp_l4_p0_col11_cout;
	wire  u_comp_l4_p0_col11_sum ;
	wire  u_comp_l4_p0_col12_cout;
	wire  u_comp_l4_p0_col12_sum ;
	wire  u_comp_l4_p0_col13_cout;
	wire  u_comp_l4_p0_col13_sum ;
	wire  u_comp_l4_p0_col14_cout;
	wire  u_comp_l4_p0_col14_sum ;
	wire  u_comp_l4_p0_col15_cout;
	wire  u_comp_l4_p0_col15_sum ;
	wire  u_comp_l4_p0_col16_cout;
	wire  u_comp_l4_p0_col16_sum ;
	wire  u_comp_l4_p0_col17_cout;
	wire  u_comp_l4_p0_col17_sum ;
	wire  u_comp_l4_p0_col18_cout;
	wire  u_comp_l4_p0_col18_sum ;
	wire  u_comp_l4_p0_col19_cout;
	wire  u_comp_l4_p0_col19_sum ;
	wire  u_comp_l4_p0_col20_cout;
	wire  u_comp_l4_p0_col20_sum ;
	wire  u_comp_l4_p0_col21_cout;
	wire  u_comp_l4_p0_col21_sum ;
	wire  u_comp_l4_p0_col22_cout;
	wire  u_comp_l4_p0_col22_sum ;
	wire  u_comp_l4_p0_col23_cout;
	wire  u_comp_l4_p0_col23_sum ;
	wire  u_comp_l4_p0_col24_cout;
	wire  u_comp_l4_p0_col24_sum ;
	wire  u_comp_l4_p0_col25_cout;
	wire  u_comp_l4_p0_col25_sum ;
	wire  u_comp_l4_p0_col26_cout;
	wire  u_comp_l4_p0_col26_sum ;
	wire  u_comp_l4_p0_col27_cout;
	wire  u_comp_l4_p0_col27_sum ;
	wire  u_comp_l4_p0_col28_cout;
	wire  u_comp_l4_p0_col28_sum ;
	wire  u_comp_l4_p0_col29_cout;
	wire  u_comp_l4_p0_col29_sum ;
	wire  u_comp_l4_p0_col30_cout;
	wire  u_comp_l4_p0_col30_sum ;
	wire  u_comp_l4_p0_col31_sum ;

	//Wire define for Inout.

	//Wire sub module connect to this module and inter module connect.
	assign p_0_0 = pp_0[0];
	
	assign p_0_1 = pp_0[1];
	
	assign p_0_2 = pp_0[2];
	
	assign p_0_3 = pp_0[3];
	
	assign p_0_4 = pp_0[4];
	
	assign p_0_5 = pp_0[5];
	
	assign p_0_6 = pp_0[6];
	
	assign p_0_7 = pp_0[7];
	
	assign p_0_8 = pp_0[8];
	
	assign p_0_9 = pp_0[9];
	
	assign p_0_10 = pp_0[10];
	
	assign p_0_11 = pp_0[11];
	
	assign p_0_12 = pp_0[12];
	
	assign p_0_13 = pp_0[13];
	
	assign p_0_14 = pp_0[14];
	
	assign p_0_15 = pp_0[15];
	
	assign p_0_16 = pp_0[16];
	
	assign p_0_17 = pp_0[17];
	
	assign p_0_18 = pp_0[18];
	
	assign p_0_19 = pp_0[19];
	
	assign p_0_20 = pp_0[20];
	
	assign p_0_21 = pp_0[21];
	
	assign p_0_22 = pp_0[22];
	
	assign p_0_23 = pp_0[23];
	
	assign p_0_24 = pp_0[24];
	
	assign p_0_25 = pp_0[25];
	
	assign p_0_26 = pp_0[26];
	
	assign p_0_27 = pp_0[27];
	
	assign p_0_28 = pp_0[28];
	
	assign p_0_29 = pp_0[29];
	
	assign p_0_30 = pp_0[30];
	
	assign p_0_31 = pp_0[31];
	
	assign p_1_0 = pp_1[0];
	
	assign p_1_1 = pp_1[1];
	
	assign p_1_2 = pp_1[2];
	
	assign p_1_3 = pp_1[3];
	
	assign p_1_4 = pp_1[4];
	
	assign p_1_5 = pp_1[5];
	
	assign p_1_6 = pp_1[6];
	
	assign p_1_7 = pp_1[7];
	
	assign p_1_8 = pp_1[8];
	
	assign p_1_9 = pp_1[9];
	
	assign p_1_10 = pp_1[10];
	
	assign p_1_11 = pp_1[11];
	
	assign p_1_12 = pp_1[12];
	
	assign p_1_13 = pp_1[13];
	
	assign p_1_14 = pp_1[14];
	
	assign p_1_15 = pp_1[15];
	
	assign p_1_16 = pp_1[16];
	
	assign p_1_17 = pp_1[17];
	
	assign p_1_18 = pp_1[18];
	
	assign p_1_19 = pp_1[19];
	
	assign p_1_20 = pp_1[20];
	
	assign p_1_21 = pp_1[21];
	
	assign p_1_22 = pp_1[22];
	
	assign p_1_23 = pp_1[23];
	
	assign p_1_24 = pp_1[24];
	
	assign p_1_25 = pp_1[25];
	
	assign p_1_26 = pp_1[26];
	
	assign p_1_27 = pp_1[27];
	
	assign p_1_28 = pp_1[28];
	
	assign p_1_29 = pp_1[29];
	
	assign p_1_30 = pp_1[30];
	
	assign p_1_31 = pp_1[31];
	
	assign p_2_0 = pp_2[0];
	
	assign p_2_1 = pp_2[1];
	
	assign p_2_2 = pp_2[2];
	
	assign p_2_3 = pp_2[3];
	
	assign p_2_4 = pp_2[4];
	
	assign p_2_5 = pp_2[5];
	
	assign p_2_6 = pp_2[6];
	
	assign p_2_7 = pp_2[7];
	
	assign p_2_8 = pp_2[8];
	
	assign p_2_9 = pp_2[9];
	
	assign p_2_10 = pp_2[10];
	
	assign p_2_11 = pp_2[11];
	
	assign p_2_12 = pp_2[12];
	
	assign p_2_13 = pp_2[13];
	
	assign p_2_14 = pp_2[14];
	
	assign p_2_15 = pp_2[15];
	
	assign p_2_16 = pp_2[16];
	
	assign p_2_17 = pp_2[17];
	
	assign p_2_18 = pp_2[18];
	
	assign p_2_19 = pp_2[19];
	
	assign p_2_20 = pp_2[20];
	
	assign p_2_21 = pp_2[21];
	
	assign p_2_22 = pp_2[22];
	
	assign p_2_23 = pp_2[23];
	
	assign p_2_24 = pp_2[24];
	
	assign p_2_25 = pp_2[25];
	
	assign p_2_26 = pp_2[26];
	
	assign p_2_27 = pp_2[27];
	
	assign p_2_28 = pp_2[28];
	
	assign p_2_29 = pp_2[29];
	
	assign p_2_30 = pp_2[30];
	
	assign p_2_31 = pp_2[31];
	
	assign p_3_0 = pp_3[0];
	
	assign p_3_1 = pp_3[1];
	
	assign p_3_2 = pp_3[2];
	
	assign p_3_3 = pp_3[3];
	
	assign p_3_4 = pp_3[4];
	
	assign p_3_5 = pp_3[5];
	
	assign p_3_6 = pp_3[6];
	
	assign p_3_7 = pp_3[7];
	
	assign p_3_8 = pp_3[8];
	
	assign p_3_9 = pp_3[9];
	
	assign p_3_10 = pp_3[10];
	
	assign p_3_11 = pp_3[11];
	
	assign p_3_12 = pp_3[12];
	
	assign p_3_13 = pp_3[13];
	
	assign p_3_14 = pp_3[14];
	
	assign p_3_15 = pp_3[15];
	
	assign p_3_16 = pp_3[16];
	
	assign p_3_17 = pp_3[17];
	
	assign p_3_18 = pp_3[18];
	
	assign p_3_19 = pp_3[19];
	
	assign p_3_20 = pp_3[20];
	
	assign p_3_21 = pp_3[21];
	
	assign p_3_22 = pp_3[22];
	
	assign p_3_23 = pp_3[23];
	
	assign p_3_24 = pp_3[24];
	
	assign p_3_25 = pp_3[25];
	
	assign p_3_26 = pp_3[26];
	
	assign p_3_27 = pp_3[27];
	
	assign p_3_28 = pp_3[28];
	
	assign p_3_29 = pp_3[29];
	
	assign p_3_30 = pp_3[30];
	
	assign p_3_31 = pp_3[31];
	
	assign p_4_0 = pp_4[0];
	
	assign p_4_1 = pp_4[1];
	
	assign p_4_2 = pp_4[2];
	
	assign p_4_3 = pp_4[3];
	
	assign p_4_4 = pp_4[4];
	
	assign p_4_5 = pp_4[5];
	
	assign p_4_6 = pp_4[6];
	
	assign p_4_7 = pp_4[7];
	
	assign p_4_8 = pp_4[8];
	
	assign p_4_9 = pp_4[9];
	
	assign p_4_10 = pp_4[10];
	
	assign p_4_11 = pp_4[11];
	
	assign p_4_12 = pp_4[12];
	
	assign p_4_13 = pp_4[13];
	
	assign p_4_14 = pp_4[14];
	
	assign p_4_15 = pp_4[15];
	
	assign p_4_16 = pp_4[16];
	
	assign p_4_17 = pp_4[17];
	
	assign p_4_18 = pp_4[18];
	
	assign p_4_19 = pp_4[19];
	
	assign p_4_20 = pp_4[20];
	
	assign p_4_21 = pp_4[21];
	
	assign p_4_22 = pp_4[22];
	
	assign p_4_23 = pp_4[23];
	
	assign p_4_24 = pp_4[24];
	
	assign p_4_25 = pp_4[25];
	
	assign p_4_26 = pp_4[26];
	
	assign p_4_27 = pp_4[27];
	
	assign p_4_28 = pp_4[28];
	
	assign p_4_29 = pp_4[29];
	
	assign p_4_30 = pp_4[30];
	
	assign p_4_31 = pp_4[31];
	
	assign p_5_0 = pp_5[0];
	
	assign p_5_1 = pp_5[1];
	
	assign p_5_2 = pp_5[2];
	
	assign p_5_3 = pp_5[3];
	
	assign p_5_4 = pp_5[4];
	
	assign p_5_5 = pp_5[5];
	
	assign p_5_6 = pp_5[6];
	
	assign p_5_7 = pp_5[7];
	
	assign p_5_8 = pp_5[8];
	
	assign p_5_9 = pp_5[9];
	
	assign p_5_10 = pp_5[10];
	
	assign p_5_11 = pp_5[11];
	
	assign p_5_12 = pp_5[12];
	
	assign p_5_13 = pp_5[13];
	
	assign p_5_14 = pp_5[14];
	
	assign p_5_15 = pp_5[15];
	
	assign p_5_16 = pp_5[16];
	
	assign p_5_17 = pp_5[17];
	
	assign p_5_18 = pp_5[18];
	
	assign p_5_19 = pp_5[19];
	
	assign p_5_20 = pp_5[20];
	
	assign p_5_21 = pp_5[21];
	
	assign p_5_22 = pp_5[22];
	
	assign p_5_23 = pp_5[23];
	
	assign p_5_24 = pp_5[24];
	
	assign p_5_25 = pp_5[25];
	
	assign p_5_26 = pp_5[26];
	
	assign p_5_27 = pp_5[27];
	
	assign p_5_28 = pp_5[28];
	
	assign p_5_29 = pp_5[29];
	
	assign p_5_30 = pp_5[30];
	
	assign p_5_31 = pp_5[31];
	
	assign p_6_0 = pp_6[0];
	
	assign p_6_1 = pp_6[1];
	
	assign p_6_2 = pp_6[2];
	
	assign p_6_3 = pp_6[3];
	
	assign p_6_4 = pp_6[4];
	
	assign p_6_5 = pp_6[5];
	
	assign p_6_6 = pp_6[6];
	
	assign p_6_7 = pp_6[7];
	
	assign p_6_8 = pp_6[8];
	
	assign p_6_9 = pp_6[9];
	
	assign p_6_10 = pp_6[10];
	
	assign p_6_11 = pp_6[11];
	
	assign p_6_12 = pp_6[12];
	
	assign p_6_13 = pp_6[13];
	
	assign p_6_14 = pp_6[14];
	
	assign p_6_15 = pp_6[15];
	
	assign p_6_16 = pp_6[16];
	
	assign p_6_17 = pp_6[17];
	
	assign p_6_18 = pp_6[18];
	
	assign p_6_19 = pp_6[19];
	
	assign p_6_20 = pp_6[20];
	
	assign p_6_21 = pp_6[21];
	
	assign p_6_22 = pp_6[22];
	
	assign p_6_23 = pp_6[23];
	
	assign p_6_24 = pp_6[24];
	
	assign p_6_25 = pp_6[25];
	
	assign p_6_26 = pp_6[26];
	
	assign p_6_27 = pp_6[27];
	
	assign p_6_28 = pp_6[28];
	
	assign p_6_29 = pp_6[29];
	
	assign p_6_30 = pp_6[30];
	
	assign p_6_31 = pp_6[31];
	
	assign p_7_0 = pp_7[0];
	
	assign p_7_1 = pp_7[1];
	
	assign p_7_2 = pp_7[2];
	
	assign p_7_3 = pp_7[3];
	
	assign p_7_4 = pp_7[4];
	
	assign p_7_5 = pp_7[5];
	
	assign p_7_6 = pp_7[6];
	
	assign p_7_7 = pp_7[7];
	
	assign p_7_8 = pp_7[8];
	
	assign p_7_9 = pp_7[9];
	
	assign p_7_10 = pp_7[10];
	
	assign p_7_11 = pp_7[11];
	
	assign p_7_12 = pp_7[12];
	
	assign p_7_13 = pp_7[13];
	
	assign p_7_14 = pp_7[14];
	
	assign p_7_15 = pp_7[15];
	
	assign p_7_16 = pp_7[16];
	
	assign p_7_17 = pp_7[17];
	
	assign p_7_18 = pp_7[18];
	
	assign p_7_19 = pp_7[19];
	
	assign p_7_20 = pp_7[20];
	
	assign p_7_21 = pp_7[21];
	
	assign p_7_22 = pp_7[22];
	
	assign p_7_23 = pp_7[23];
	
	assign p_7_24 = pp_7[24];
	
	assign p_7_25 = pp_7[25];
	
	assign p_7_26 = pp_7[26];
	
	assign p_7_27 = pp_7[27];
	
	assign p_7_28 = pp_7[28];
	
	assign p_7_29 = pp_7[29];
	
	assign p_7_30 = pp_7[30];
	
	assign p_7_31 = pp_7[31];
	
	assign p_8_0 = pp_8[0];
	
	assign p_8_1 = pp_8[1];
	
	assign p_8_2 = pp_8[2];
	
	assign p_8_3 = pp_8[3];
	
	assign p_8_4 = pp_8[4];
	
	assign p_8_5 = pp_8[5];
	
	assign p_8_6 = pp_8[6];
	
	assign p_8_7 = pp_8[7];
	
	assign p_8_8 = pp_8[8];
	
	assign p_8_9 = pp_8[9];
	
	assign p_8_10 = pp_8[10];
	
	assign p_8_11 = pp_8[11];
	
	assign p_8_12 = pp_8[12];
	
	assign p_8_13 = pp_8[13];
	
	assign p_8_14 = pp_8[14];
	
	assign p_8_15 = pp_8[15];
	
	assign p_8_16 = pp_8[16];
	
	assign p_8_17 = pp_8[17];
	
	assign p_8_18 = pp_8[18];
	
	assign p_8_19 = pp_8[19];
	
	assign p_8_20 = pp_8[20];
	
	assign p_8_21 = pp_8[21];
	
	assign p_8_22 = pp_8[22];
	
	assign p_8_23 = pp_8[23];
	
	assign p_8_24 = pp_8[24];
	
	assign p_8_25 = pp_8[25];
	
	assign p_8_26 = pp_8[26];
	
	assign p_8_27 = pp_8[27];
	
	assign p_8_28 = pp_8[28];
	
	assign p_8_29 = pp_8[29];
	
	assign p_8_30 = pp_8[30];
	
	assign p_8_31 = pp_8[31];
	
	assign p_9_0 = pp_9[0];
	
	assign p_9_1 = pp_9[1];
	
	assign p_9_2 = pp_9[2];
	
	assign p_9_3 = pp_9[3];
	
	assign p_9_4 = pp_9[4];
	
	assign p_9_5 = pp_9[5];
	
	assign p_9_6 = pp_9[6];
	
	assign p_9_7 = pp_9[7];
	
	assign p_9_8 = pp_9[8];
	
	assign p_9_9 = pp_9[9];
	
	assign p_9_10 = pp_9[10];
	
	assign p_9_11 = pp_9[11];
	
	assign p_9_12 = pp_9[12];
	
	assign p_9_13 = pp_9[13];
	
	assign p_9_14 = pp_9[14];
	
	assign p_9_15 = pp_9[15];
	
	assign p_9_16 = pp_9[16];
	
	assign p_9_17 = pp_9[17];
	
	assign p_9_18 = pp_9[18];
	
	assign p_9_19 = pp_9[19];
	
	assign p_9_20 = pp_9[20];
	
	assign p_9_21 = pp_9[21];
	
	assign p_9_22 = pp_9[22];
	
	assign p_9_23 = pp_9[23];
	
	assign p_9_24 = pp_9[24];
	
	assign p_9_25 = pp_9[25];
	
	assign p_9_26 = pp_9[26];
	
	assign p_9_27 = pp_9[27];
	
	assign p_9_28 = pp_9[28];
	
	assign p_9_29 = pp_9[29];
	
	assign p_9_30 = pp_9[30];
	
	assign p_9_31 = pp_9[31];
	
	assign ps_0 = {comp_l4_p0_col31_sum, comp_l4_p0_col30_sum, comp_l4_p0_col29_sum, comp_l4_p0_col28_sum, comp_l4_p0_col27_sum, comp_l4_p0_col26_sum, comp_l4_p0_col25_sum, comp_l4_p0_col24_sum, comp_l4_p0_col23_sum, comp_l4_p0_col22_sum, comp_l4_p0_col21_sum, comp_l4_p0_col20_sum, comp_l4_p0_col19_sum, comp_l4_p0_col18_sum, comp_l4_p0_col17_sum, comp_l4_p0_col16_sum, comp_l4_p0_col15_sum, comp_l4_p0_col14_sum, comp_l4_p0_col13_sum, comp_l4_p0_col12_sum, comp_l4_p0_col11_sum, comp_l4_p0_col10_sum, comp_l4_p0_col9_sum, comp_l4_p0_col8_sum, comp_l4_p0_col7_sum, comp_l4_p0_col6_sum, comp_l4_p0_col5_sum, comp_l4_p0_col4_sum, comp_l4_p0_col3_sum, comp_l4_p0_col2_sum, comp_l4_p0_col1_sum, comp_l4_p0_col0_sum};
	
	assign ps_1 = {comp_l4_p0_col30_cout, comp_l4_p0_col29_cout, comp_l4_p0_col28_cout, comp_l4_p0_col27_cout, comp_l4_p0_col26_cout, comp_l4_p0_col25_cout, comp_l4_p0_col24_cout, comp_l4_p0_col23_cout, comp_l4_p0_col22_cout, comp_l4_p0_col21_cout, comp_l4_p0_col20_cout, comp_l4_p0_col19_cout, comp_l4_p0_col18_cout, comp_l4_p0_col17_cout, comp_l4_p0_col16_cout, comp_l4_p0_col15_cout, comp_l4_p0_col14_cout, comp_l4_p0_col13_cout, comp_l4_p0_col12_cout, comp_l4_p0_col11_cout, comp_l4_p0_col10_cout, comp_l4_p0_col9_cout, comp_l4_p0_col8_cout, comp_l4_p0_col7_cout, comp_l4_p0_col6_cout, comp_l4_p0_col5_cout, comp_l4_p0_col4_cout, comp_l4_p0_col3_cout, comp_l4_p0_col2_cout, comp_l4_p0_col1_cout, comp_l4_p0_col0_cout, comp_pad_l4_p0};
	
	assign comp_l0_p0_col0_cout = u_comp_l0_p0_col0_cout;
	
	assign comp_l0_p0_col0_sum = u_comp_l0_p0_col0_sum;
	
	assign comp_l0_p0_col1_cout = u_comp_l0_p0_col1_cout;
	
	assign comp_l0_p0_col1_sum = u_comp_l0_p0_col1_sum;
	
	assign comp_l0_p0_col2_cout = u_comp_l0_p0_col2_cout;
	
	assign comp_l0_p0_col2_sum = u_comp_l0_p0_col2_sum;
	
	assign comp_l0_p0_col3_cout = u_comp_l0_p0_col3_cout;
	
	assign comp_l0_p0_col3_sum = u_comp_l0_p0_col3_sum;
	
	assign comp_l0_p0_col4_cout = u_comp_l0_p0_col4_cout;
	
	assign comp_l0_p0_col4_sum = u_comp_l0_p0_col4_sum;
	
	assign comp_l0_p0_col5_cout = u_comp_l0_p0_col5_cout;
	
	assign comp_l0_p0_col5_sum = u_comp_l0_p0_col5_sum;
	
	assign comp_l0_p0_col6_cout = u_comp_l0_p0_col6_cout;
	
	assign comp_l0_p0_col6_sum = u_comp_l0_p0_col6_sum;
	
	assign comp_l0_p0_col7_cout = u_comp_l0_p0_col7_cout;
	
	assign comp_l0_p0_col7_sum = u_comp_l0_p0_col7_sum;
	
	assign comp_l0_p0_col8_cout = u_comp_l0_p0_col8_cout;
	
	assign comp_l0_p0_col8_sum = u_comp_l0_p0_col8_sum;
	
	assign comp_l0_p0_col9_cout = u_comp_l0_p0_col9_cout;
	
	assign comp_l0_p0_col9_sum = u_comp_l0_p0_col9_sum;
	
	assign comp_l0_p0_col10_cout = u_comp_l0_p0_col10_cout;
	
	assign comp_l0_p0_col10_sum = u_comp_l0_p0_col10_sum;
	
	assign comp_l0_p0_col11_cout = u_comp_l0_p0_col11_cout;
	
	assign comp_l0_p0_col11_sum = u_comp_l0_p0_col11_sum;
	
	assign comp_l0_p0_col12_cout = u_comp_l0_p0_col12_cout;
	
	assign comp_l0_p0_col12_sum = u_comp_l0_p0_col12_sum;
	
	assign comp_l0_p0_col13_cout = u_comp_l0_p0_col13_cout;
	
	assign comp_l0_p0_col13_sum = u_comp_l0_p0_col13_sum;
	
	assign comp_l0_p0_col14_cout = u_comp_l0_p0_col14_cout;
	
	assign comp_l0_p0_col14_sum = u_comp_l0_p0_col14_sum;
	
	assign comp_l0_p0_col15_cout = u_comp_l0_p0_col15_cout;
	
	assign comp_l0_p0_col15_sum = u_comp_l0_p0_col15_sum;
	
	assign comp_l0_p0_col16_cout = u_comp_l0_p0_col16_cout;
	
	assign comp_l0_p0_col16_sum = u_comp_l0_p0_col16_sum;
	
	assign comp_l0_p0_col17_cout = u_comp_l0_p0_col17_cout;
	
	assign comp_l0_p0_col17_sum = u_comp_l0_p0_col17_sum;
	
	assign comp_l0_p0_col18_cout = u_comp_l0_p0_col18_cout;
	
	assign comp_l0_p0_col18_sum = u_comp_l0_p0_col18_sum;
	
	assign comp_l0_p0_col19_cout = u_comp_l0_p0_col19_cout;
	
	assign comp_l0_p0_col19_sum = u_comp_l0_p0_col19_sum;
	
	assign comp_l0_p0_col20_cout = u_comp_l0_p0_col20_cout;
	
	assign comp_l0_p0_col20_sum = u_comp_l0_p0_col20_sum;
	
	assign comp_l0_p0_col21_cout = u_comp_l0_p0_col21_cout;
	
	assign comp_l0_p0_col21_sum = u_comp_l0_p0_col21_sum;
	
	assign comp_l0_p0_col22_cout = u_comp_l0_p0_col22_cout;
	
	assign comp_l0_p0_col22_sum = u_comp_l0_p0_col22_sum;
	
	assign comp_l0_p0_col23_cout = u_comp_l0_p0_col23_cout;
	
	assign comp_l0_p0_col23_sum = u_comp_l0_p0_col23_sum;
	
	assign comp_l0_p0_col24_cout = u_comp_l0_p0_col24_cout;
	
	assign comp_l0_p0_col24_sum = u_comp_l0_p0_col24_sum;
	
	assign comp_l0_p0_col25_cout = u_comp_l0_p0_col25_cout;
	
	assign comp_l0_p0_col25_sum = u_comp_l0_p0_col25_sum;
	
	assign comp_l0_p0_col26_cout = u_comp_l0_p0_col26_cout;
	
	assign comp_l0_p0_col26_sum = u_comp_l0_p0_col26_sum;
	
	assign comp_l0_p0_col27_cout = u_comp_l0_p0_col27_cout;
	
	assign comp_l0_p0_col27_sum = u_comp_l0_p0_col27_sum;
	
	assign comp_l0_p0_col28_cout = u_comp_l0_p0_col28_cout;
	
	assign comp_l0_p0_col28_sum = u_comp_l0_p0_col28_sum;
	
	assign comp_l0_p0_col29_cout = u_comp_l0_p0_col29_cout;
	
	assign comp_l0_p0_col29_sum = u_comp_l0_p0_col29_sum;
	
	assign comp_l0_p0_col30_cout = u_comp_l0_p0_col30_cout;
	
	assign comp_l0_p0_col30_sum = u_comp_l0_p0_col30_sum;
	
	assign comp_l0_p0_col31_sum = u_comp_l0_p0_col31_sum;
	
	assign comp_pad_l0_p0 = 1'b0;
	
	assign comp_l0_p1_col0_cout = u_comp_l0_p1_col0_cout;
	
	assign comp_l0_p1_col0_sum = u_comp_l0_p1_col0_sum;
	
	assign comp_l0_p1_col1_cout = u_comp_l0_p1_col1_cout;
	
	assign comp_l0_p1_col1_sum = u_comp_l0_p1_col1_sum;
	
	assign comp_l0_p1_col2_cout = u_comp_l0_p1_col2_cout;
	
	assign comp_l0_p1_col2_sum = u_comp_l0_p1_col2_sum;
	
	assign comp_l0_p1_col3_cout = u_comp_l0_p1_col3_cout;
	
	assign comp_l0_p1_col3_sum = u_comp_l0_p1_col3_sum;
	
	assign comp_l0_p1_col4_cout = u_comp_l0_p1_col4_cout;
	
	assign comp_l0_p1_col4_sum = u_comp_l0_p1_col4_sum;
	
	assign comp_l0_p1_col5_cout = u_comp_l0_p1_col5_cout;
	
	assign comp_l0_p1_col5_sum = u_comp_l0_p1_col5_sum;
	
	assign comp_l0_p1_col6_cout = u_comp_l0_p1_col6_cout;
	
	assign comp_l0_p1_col6_sum = u_comp_l0_p1_col6_sum;
	
	assign comp_l0_p1_col7_cout = u_comp_l0_p1_col7_cout;
	
	assign comp_l0_p1_col7_sum = u_comp_l0_p1_col7_sum;
	
	assign comp_l0_p1_col8_cout = u_comp_l0_p1_col8_cout;
	
	assign comp_l0_p1_col8_sum = u_comp_l0_p1_col8_sum;
	
	assign comp_l0_p1_col9_cout = u_comp_l0_p1_col9_cout;
	
	assign comp_l0_p1_col9_sum = u_comp_l0_p1_col9_sum;
	
	assign comp_l0_p1_col10_cout = u_comp_l0_p1_col10_cout;
	
	assign comp_l0_p1_col10_sum = u_comp_l0_p1_col10_sum;
	
	assign comp_l0_p1_col11_cout = u_comp_l0_p1_col11_cout;
	
	assign comp_l0_p1_col11_sum = u_comp_l0_p1_col11_sum;
	
	assign comp_l0_p1_col12_cout = u_comp_l0_p1_col12_cout;
	
	assign comp_l0_p1_col12_sum = u_comp_l0_p1_col12_sum;
	
	assign comp_l0_p1_col13_cout = u_comp_l0_p1_col13_cout;
	
	assign comp_l0_p1_col13_sum = u_comp_l0_p1_col13_sum;
	
	assign comp_l0_p1_col14_cout = u_comp_l0_p1_col14_cout;
	
	assign comp_l0_p1_col14_sum = u_comp_l0_p1_col14_sum;
	
	assign comp_l0_p1_col15_cout = u_comp_l0_p1_col15_cout;
	
	assign comp_l0_p1_col15_sum = u_comp_l0_p1_col15_sum;
	
	assign comp_l0_p1_col16_cout = u_comp_l0_p1_col16_cout;
	
	assign comp_l0_p1_col16_sum = u_comp_l0_p1_col16_sum;
	
	assign comp_l0_p1_col17_cout = u_comp_l0_p1_col17_cout;
	
	assign comp_l0_p1_col17_sum = u_comp_l0_p1_col17_sum;
	
	assign comp_l0_p1_col18_cout = u_comp_l0_p1_col18_cout;
	
	assign comp_l0_p1_col18_sum = u_comp_l0_p1_col18_sum;
	
	assign comp_l0_p1_col19_cout = u_comp_l0_p1_col19_cout;
	
	assign comp_l0_p1_col19_sum = u_comp_l0_p1_col19_sum;
	
	assign comp_l0_p1_col20_cout = u_comp_l0_p1_col20_cout;
	
	assign comp_l0_p1_col20_sum = u_comp_l0_p1_col20_sum;
	
	assign comp_l0_p1_col21_cout = u_comp_l0_p1_col21_cout;
	
	assign comp_l0_p1_col21_sum = u_comp_l0_p1_col21_sum;
	
	assign comp_l0_p1_col22_cout = u_comp_l0_p1_col22_cout;
	
	assign comp_l0_p1_col22_sum = u_comp_l0_p1_col22_sum;
	
	assign comp_l0_p1_col23_cout = u_comp_l0_p1_col23_cout;
	
	assign comp_l0_p1_col23_sum = u_comp_l0_p1_col23_sum;
	
	assign comp_l0_p1_col24_cout = u_comp_l0_p1_col24_cout;
	
	assign comp_l0_p1_col24_sum = u_comp_l0_p1_col24_sum;
	
	assign comp_l0_p1_col25_cout = u_comp_l0_p1_col25_cout;
	
	assign comp_l0_p1_col25_sum = u_comp_l0_p1_col25_sum;
	
	assign comp_l0_p1_col26_cout = u_comp_l0_p1_col26_cout;
	
	assign comp_l0_p1_col26_sum = u_comp_l0_p1_col26_sum;
	
	assign comp_l0_p1_col27_cout = u_comp_l0_p1_col27_cout;
	
	assign comp_l0_p1_col27_sum = u_comp_l0_p1_col27_sum;
	
	assign comp_l0_p1_col28_cout = u_comp_l0_p1_col28_cout;
	
	assign comp_l0_p1_col28_sum = u_comp_l0_p1_col28_sum;
	
	assign comp_l0_p1_col29_cout = u_comp_l0_p1_col29_cout;
	
	assign comp_l0_p1_col29_sum = u_comp_l0_p1_col29_sum;
	
	assign comp_l0_p1_col30_cout = u_comp_l0_p1_col30_cout;
	
	assign comp_l0_p1_col30_sum = u_comp_l0_p1_col30_sum;
	
	assign comp_l0_p1_col31_sum = u_comp_l0_p1_col31_sum;
	
	assign comp_pad_l0_p1 = 1'b0;
	
	assign comp_l0_p2_col0_cout = u_comp_l0_p2_col0_cout;
	
	assign comp_l0_p2_col0_sum = u_comp_l0_p2_col0_sum;
	
	assign comp_l0_p2_col1_cout = u_comp_l0_p2_col1_cout;
	
	assign comp_l0_p2_col1_sum = u_comp_l0_p2_col1_sum;
	
	assign comp_l0_p2_col2_cout = u_comp_l0_p2_col2_cout;
	
	assign comp_l0_p2_col2_sum = u_comp_l0_p2_col2_sum;
	
	assign comp_l0_p2_col3_cout = u_comp_l0_p2_col3_cout;
	
	assign comp_l0_p2_col3_sum = u_comp_l0_p2_col3_sum;
	
	assign comp_l0_p2_col4_cout = u_comp_l0_p2_col4_cout;
	
	assign comp_l0_p2_col4_sum = u_comp_l0_p2_col4_sum;
	
	assign comp_l0_p2_col5_cout = u_comp_l0_p2_col5_cout;
	
	assign comp_l0_p2_col5_sum = u_comp_l0_p2_col5_sum;
	
	assign comp_l0_p2_col6_cout = u_comp_l0_p2_col6_cout;
	
	assign comp_l0_p2_col6_sum = u_comp_l0_p2_col6_sum;
	
	assign comp_l0_p2_col7_cout = u_comp_l0_p2_col7_cout;
	
	assign comp_l0_p2_col7_sum = u_comp_l0_p2_col7_sum;
	
	assign comp_l0_p2_col8_cout = u_comp_l0_p2_col8_cout;
	
	assign comp_l0_p2_col8_sum = u_comp_l0_p2_col8_sum;
	
	assign comp_l0_p2_col9_cout = u_comp_l0_p2_col9_cout;
	
	assign comp_l0_p2_col9_sum = u_comp_l0_p2_col9_sum;
	
	assign comp_l0_p2_col10_cout = u_comp_l0_p2_col10_cout;
	
	assign comp_l0_p2_col10_sum = u_comp_l0_p2_col10_sum;
	
	assign comp_l0_p2_col11_cout = u_comp_l0_p2_col11_cout;
	
	assign comp_l0_p2_col11_sum = u_comp_l0_p2_col11_sum;
	
	assign comp_l0_p2_col12_cout = u_comp_l0_p2_col12_cout;
	
	assign comp_l0_p2_col12_sum = u_comp_l0_p2_col12_sum;
	
	assign comp_l0_p2_col13_cout = u_comp_l0_p2_col13_cout;
	
	assign comp_l0_p2_col13_sum = u_comp_l0_p2_col13_sum;
	
	assign comp_l0_p2_col14_cout = u_comp_l0_p2_col14_cout;
	
	assign comp_l0_p2_col14_sum = u_comp_l0_p2_col14_sum;
	
	assign comp_l0_p2_col15_cout = u_comp_l0_p2_col15_cout;
	
	assign comp_l0_p2_col15_sum = u_comp_l0_p2_col15_sum;
	
	assign comp_l0_p2_col16_cout = u_comp_l0_p2_col16_cout;
	
	assign comp_l0_p2_col16_sum = u_comp_l0_p2_col16_sum;
	
	assign comp_l0_p2_col17_cout = u_comp_l0_p2_col17_cout;
	
	assign comp_l0_p2_col17_sum = u_comp_l0_p2_col17_sum;
	
	assign comp_l0_p2_col18_cout = u_comp_l0_p2_col18_cout;
	
	assign comp_l0_p2_col18_sum = u_comp_l0_p2_col18_sum;
	
	assign comp_l0_p2_col19_cout = u_comp_l0_p2_col19_cout;
	
	assign comp_l0_p2_col19_sum = u_comp_l0_p2_col19_sum;
	
	assign comp_l0_p2_col20_cout = u_comp_l0_p2_col20_cout;
	
	assign comp_l0_p2_col20_sum = u_comp_l0_p2_col20_sum;
	
	assign comp_l0_p2_col21_cout = u_comp_l0_p2_col21_cout;
	
	assign comp_l0_p2_col21_sum = u_comp_l0_p2_col21_sum;
	
	assign comp_l0_p2_col22_cout = u_comp_l0_p2_col22_cout;
	
	assign comp_l0_p2_col22_sum = u_comp_l0_p2_col22_sum;
	
	assign comp_l0_p2_col23_cout = u_comp_l0_p2_col23_cout;
	
	assign comp_l0_p2_col23_sum = u_comp_l0_p2_col23_sum;
	
	assign comp_l0_p2_col24_cout = u_comp_l0_p2_col24_cout;
	
	assign comp_l0_p2_col24_sum = u_comp_l0_p2_col24_sum;
	
	assign comp_l0_p2_col25_cout = u_comp_l0_p2_col25_cout;
	
	assign comp_l0_p2_col25_sum = u_comp_l0_p2_col25_sum;
	
	assign comp_l0_p2_col26_cout = u_comp_l0_p2_col26_cout;
	
	assign comp_l0_p2_col26_sum = u_comp_l0_p2_col26_sum;
	
	assign comp_l0_p2_col27_cout = u_comp_l0_p2_col27_cout;
	
	assign comp_l0_p2_col27_sum = u_comp_l0_p2_col27_sum;
	
	assign comp_l0_p2_col28_cout = u_comp_l0_p2_col28_cout;
	
	assign comp_l0_p2_col28_sum = u_comp_l0_p2_col28_sum;
	
	assign comp_l0_p2_col29_cout = u_comp_l0_p2_col29_cout;
	
	assign comp_l0_p2_col29_sum = u_comp_l0_p2_col29_sum;
	
	assign comp_l0_p2_col30_cout = u_comp_l0_p2_col30_cout;
	
	assign comp_l0_p2_col30_sum = u_comp_l0_p2_col30_sum;
	
	assign comp_l0_p2_col31_sum = u_comp_l0_p2_col31_sum;
	
	assign comp_pad_l0_p2 = 1'b0;
	
	assign comp_l1_p0_col0_cout = u_comp_l1_p0_col0_cout;
	
	assign comp_l1_p0_col0_sum = u_comp_l1_p0_col0_sum;
	
	assign comp_l1_p0_col1_cout = u_comp_l1_p0_col1_cout;
	
	assign comp_l1_p0_col1_sum = u_comp_l1_p0_col1_sum;
	
	assign comp_l1_p0_col2_cout = u_comp_l1_p0_col2_cout;
	
	assign comp_l1_p0_col2_sum = u_comp_l1_p0_col2_sum;
	
	assign comp_l1_p0_col3_cout = u_comp_l1_p0_col3_cout;
	
	assign comp_l1_p0_col3_sum = u_comp_l1_p0_col3_sum;
	
	assign comp_l1_p0_col4_cout = u_comp_l1_p0_col4_cout;
	
	assign comp_l1_p0_col4_sum = u_comp_l1_p0_col4_sum;
	
	assign comp_l1_p0_col5_cout = u_comp_l1_p0_col5_cout;
	
	assign comp_l1_p0_col5_sum = u_comp_l1_p0_col5_sum;
	
	assign comp_l1_p0_col6_cout = u_comp_l1_p0_col6_cout;
	
	assign comp_l1_p0_col6_sum = u_comp_l1_p0_col6_sum;
	
	assign comp_l1_p0_col7_cout = u_comp_l1_p0_col7_cout;
	
	assign comp_l1_p0_col7_sum = u_comp_l1_p0_col7_sum;
	
	assign comp_l1_p0_col8_cout = u_comp_l1_p0_col8_cout;
	
	assign comp_l1_p0_col8_sum = u_comp_l1_p0_col8_sum;
	
	assign comp_l1_p0_col9_cout = u_comp_l1_p0_col9_cout;
	
	assign comp_l1_p0_col9_sum = u_comp_l1_p0_col9_sum;
	
	assign comp_l1_p0_col10_cout = u_comp_l1_p0_col10_cout;
	
	assign comp_l1_p0_col10_sum = u_comp_l1_p0_col10_sum;
	
	assign comp_l1_p0_col11_cout = u_comp_l1_p0_col11_cout;
	
	assign comp_l1_p0_col11_sum = u_comp_l1_p0_col11_sum;
	
	assign comp_l1_p0_col12_cout = u_comp_l1_p0_col12_cout;
	
	assign comp_l1_p0_col12_sum = u_comp_l1_p0_col12_sum;
	
	assign comp_l1_p0_col13_cout = u_comp_l1_p0_col13_cout;
	
	assign comp_l1_p0_col13_sum = u_comp_l1_p0_col13_sum;
	
	assign comp_l1_p0_col14_cout = u_comp_l1_p0_col14_cout;
	
	assign comp_l1_p0_col14_sum = u_comp_l1_p0_col14_sum;
	
	assign comp_l1_p0_col15_cout = u_comp_l1_p0_col15_cout;
	
	assign comp_l1_p0_col15_sum = u_comp_l1_p0_col15_sum;
	
	assign comp_l1_p0_col16_cout = u_comp_l1_p0_col16_cout;
	
	assign comp_l1_p0_col16_sum = u_comp_l1_p0_col16_sum;
	
	assign comp_l1_p0_col17_cout = u_comp_l1_p0_col17_cout;
	
	assign comp_l1_p0_col17_sum = u_comp_l1_p0_col17_sum;
	
	assign comp_l1_p0_col18_cout = u_comp_l1_p0_col18_cout;
	
	assign comp_l1_p0_col18_sum = u_comp_l1_p0_col18_sum;
	
	assign comp_l1_p0_col19_cout = u_comp_l1_p0_col19_cout;
	
	assign comp_l1_p0_col19_sum = u_comp_l1_p0_col19_sum;
	
	assign comp_l1_p0_col20_cout = u_comp_l1_p0_col20_cout;
	
	assign comp_l1_p0_col20_sum = u_comp_l1_p0_col20_sum;
	
	assign comp_l1_p0_col21_cout = u_comp_l1_p0_col21_cout;
	
	assign comp_l1_p0_col21_sum = u_comp_l1_p0_col21_sum;
	
	assign comp_l1_p0_col22_cout = u_comp_l1_p0_col22_cout;
	
	assign comp_l1_p0_col22_sum = u_comp_l1_p0_col22_sum;
	
	assign comp_l1_p0_col23_cout = u_comp_l1_p0_col23_cout;
	
	assign comp_l1_p0_col23_sum = u_comp_l1_p0_col23_sum;
	
	assign comp_l1_p0_col24_cout = u_comp_l1_p0_col24_cout;
	
	assign comp_l1_p0_col24_sum = u_comp_l1_p0_col24_sum;
	
	assign comp_l1_p0_col25_cout = u_comp_l1_p0_col25_cout;
	
	assign comp_l1_p0_col25_sum = u_comp_l1_p0_col25_sum;
	
	assign comp_l1_p0_col26_cout = u_comp_l1_p0_col26_cout;
	
	assign comp_l1_p0_col26_sum = u_comp_l1_p0_col26_sum;
	
	assign comp_l1_p0_col27_cout = u_comp_l1_p0_col27_cout;
	
	assign comp_l1_p0_col27_sum = u_comp_l1_p0_col27_sum;
	
	assign comp_l1_p0_col28_cout = u_comp_l1_p0_col28_cout;
	
	assign comp_l1_p0_col28_sum = u_comp_l1_p0_col28_sum;
	
	assign comp_l1_p0_col29_cout = u_comp_l1_p0_col29_cout;
	
	assign comp_l1_p0_col29_sum = u_comp_l1_p0_col29_sum;
	
	assign comp_l1_p0_col30_cout = u_comp_l1_p0_col30_cout;
	
	assign comp_l1_p0_col30_sum = u_comp_l1_p0_col30_sum;
	
	assign comp_l1_p0_col31_sum = u_comp_l1_p0_col31_sum;
	
	assign comp_pad_l1_p0 = 1'b0;
	
	assign comp_l1_p1_col0_cout = u_comp_l1_p1_col0_cout;
	
	assign comp_l1_p1_col0_sum = u_comp_l1_p1_col0_sum;
	
	assign comp_l1_p1_col1_cout = u_comp_l1_p1_col1_cout;
	
	assign comp_l1_p1_col1_sum = u_comp_l1_p1_col1_sum;
	
	assign comp_l1_p1_col2_cout = u_comp_l1_p1_col2_cout;
	
	assign comp_l1_p1_col2_sum = u_comp_l1_p1_col2_sum;
	
	assign comp_l1_p1_col3_cout = u_comp_l1_p1_col3_cout;
	
	assign comp_l1_p1_col3_sum = u_comp_l1_p1_col3_sum;
	
	assign comp_l1_p1_col4_cout = u_comp_l1_p1_col4_cout;
	
	assign comp_l1_p1_col4_sum = u_comp_l1_p1_col4_sum;
	
	assign comp_l1_p1_col5_cout = u_comp_l1_p1_col5_cout;
	
	assign comp_l1_p1_col5_sum = u_comp_l1_p1_col5_sum;
	
	assign comp_l1_p1_col6_cout = u_comp_l1_p1_col6_cout;
	
	assign comp_l1_p1_col6_sum = u_comp_l1_p1_col6_sum;
	
	assign comp_l1_p1_col7_cout = u_comp_l1_p1_col7_cout;
	
	assign comp_l1_p1_col7_sum = u_comp_l1_p1_col7_sum;
	
	assign comp_l1_p1_col8_cout = u_comp_l1_p1_col8_cout;
	
	assign comp_l1_p1_col8_sum = u_comp_l1_p1_col8_sum;
	
	assign comp_l1_p1_col9_cout = u_comp_l1_p1_col9_cout;
	
	assign comp_l1_p1_col9_sum = u_comp_l1_p1_col9_sum;
	
	assign comp_l1_p1_col10_cout = u_comp_l1_p1_col10_cout;
	
	assign comp_l1_p1_col10_sum = u_comp_l1_p1_col10_sum;
	
	assign comp_l1_p1_col11_cout = u_comp_l1_p1_col11_cout;
	
	assign comp_l1_p1_col11_sum = u_comp_l1_p1_col11_sum;
	
	assign comp_l1_p1_col12_cout = u_comp_l1_p1_col12_cout;
	
	assign comp_l1_p1_col12_sum = u_comp_l1_p1_col12_sum;
	
	assign comp_l1_p1_col13_cout = u_comp_l1_p1_col13_cout;
	
	assign comp_l1_p1_col13_sum = u_comp_l1_p1_col13_sum;
	
	assign comp_l1_p1_col14_cout = u_comp_l1_p1_col14_cout;
	
	assign comp_l1_p1_col14_sum = u_comp_l1_p1_col14_sum;
	
	assign comp_l1_p1_col15_cout = u_comp_l1_p1_col15_cout;
	
	assign comp_l1_p1_col15_sum = u_comp_l1_p1_col15_sum;
	
	assign comp_l1_p1_col16_cout = u_comp_l1_p1_col16_cout;
	
	assign comp_l1_p1_col16_sum = u_comp_l1_p1_col16_sum;
	
	assign comp_l1_p1_col17_cout = u_comp_l1_p1_col17_cout;
	
	assign comp_l1_p1_col17_sum = u_comp_l1_p1_col17_sum;
	
	assign comp_l1_p1_col18_cout = u_comp_l1_p1_col18_cout;
	
	assign comp_l1_p1_col18_sum = u_comp_l1_p1_col18_sum;
	
	assign comp_l1_p1_col19_cout = u_comp_l1_p1_col19_cout;
	
	assign comp_l1_p1_col19_sum = u_comp_l1_p1_col19_sum;
	
	assign comp_l1_p1_col20_cout = u_comp_l1_p1_col20_cout;
	
	assign comp_l1_p1_col20_sum = u_comp_l1_p1_col20_sum;
	
	assign comp_l1_p1_col21_cout = u_comp_l1_p1_col21_cout;
	
	assign comp_l1_p1_col21_sum = u_comp_l1_p1_col21_sum;
	
	assign comp_l1_p1_col22_cout = u_comp_l1_p1_col22_cout;
	
	assign comp_l1_p1_col22_sum = u_comp_l1_p1_col22_sum;
	
	assign comp_l1_p1_col23_cout = u_comp_l1_p1_col23_cout;
	
	assign comp_l1_p1_col23_sum = u_comp_l1_p1_col23_sum;
	
	assign comp_l1_p1_col24_cout = u_comp_l1_p1_col24_cout;
	
	assign comp_l1_p1_col24_sum = u_comp_l1_p1_col24_sum;
	
	assign comp_l1_p1_col25_cout = u_comp_l1_p1_col25_cout;
	
	assign comp_l1_p1_col25_sum = u_comp_l1_p1_col25_sum;
	
	assign comp_l1_p1_col26_cout = u_comp_l1_p1_col26_cout;
	
	assign comp_l1_p1_col26_sum = u_comp_l1_p1_col26_sum;
	
	assign comp_l1_p1_col27_cout = u_comp_l1_p1_col27_cout;
	
	assign comp_l1_p1_col27_sum = u_comp_l1_p1_col27_sum;
	
	assign comp_l1_p1_col28_cout = u_comp_l1_p1_col28_cout;
	
	assign comp_l1_p1_col28_sum = u_comp_l1_p1_col28_sum;
	
	assign comp_l1_p1_col29_cout = u_comp_l1_p1_col29_cout;
	
	assign comp_l1_p1_col29_sum = u_comp_l1_p1_col29_sum;
	
	assign comp_l1_p1_col30_cout = u_comp_l1_p1_col30_cout;
	
	assign comp_l1_p1_col30_sum = u_comp_l1_p1_col30_sum;
	
	assign comp_l1_p1_col31_sum = u_comp_l1_p1_col31_sum;
	
	assign comp_pad_l1_p1 = 1'b0;
	
	assign comp_l2_p0_col0_cout = u_comp_l2_p0_col0_cout;
	
	assign comp_l2_p0_col0_sum = u_comp_l2_p0_col0_sum;
	
	assign comp_l2_p0_col1_cout = u_comp_l2_p0_col1_cout;
	
	assign comp_l2_p0_col1_sum = u_comp_l2_p0_col1_sum;
	
	assign comp_l2_p0_col2_cout = u_comp_l2_p0_col2_cout;
	
	assign comp_l2_p0_col2_sum = u_comp_l2_p0_col2_sum;
	
	assign comp_l2_p0_col3_cout = u_comp_l2_p0_col3_cout;
	
	assign comp_l2_p0_col3_sum = u_comp_l2_p0_col3_sum;
	
	assign comp_l2_p0_col4_cout = u_comp_l2_p0_col4_cout;
	
	assign comp_l2_p0_col4_sum = u_comp_l2_p0_col4_sum;
	
	assign comp_l2_p0_col5_cout = u_comp_l2_p0_col5_cout;
	
	assign comp_l2_p0_col5_sum = u_comp_l2_p0_col5_sum;
	
	assign comp_l2_p0_col6_cout = u_comp_l2_p0_col6_cout;
	
	assign comp_l2_p0_col6_sum = u_comp_l2_p0_col6_sum;
	
	assign comp_l2_p0_col7_cout = u_comp_l2_p0_col7_cout;
	
	assign comp_l2_p0_col7_sum = u_comp_l2_p0_col7_sum;
	
	assign comp_l2_p0_col8_cout = u_comp_l2_p0_col8_cout;
	
	assign comp_l2_p0_col8_sum = u_comp_l2_p0_col8_sum;
	
	assign comp_l2_p0_col9_cout = u_comp_l2_p0_col9_cout;
	
	assign comp_l2_p0_col9_sum = u_comp_l2_p0_col9_sum;
	
	assign comp_l2_p0_col10_cout = u_comp_l2_p0_col10_cout;
	
	assign comp_l2_p0_col10_sum = u_comp_l2_p0_col10_sum;
	
	assign comp_l2_p0_col11_cout = u_comp_l2_p0_col11_cout;
	
	assign comp_l2_p0_col11_sum = u_comp_l2_p0_col11_sum;
	
	assign comp_l2_p0_col12_cout = u_comp_l2_p0_col12_cout;
	
	assign comp_l2_p0_col12_sum = u_comp_l2_p0_col12_sum;
	
	assign comp_l2_p0_col13_cout = u_comp_l2_p0_col13_cout;
	
	assign comp_l2_p0_col13_sum = u_comp_l2_p0_col13_sum;
	
	assign comp_l2_p0_col14_cout = u_comp_l2_p0_col14_cout;
	
	assign comp_l2_p0_col14_sum = u_comp_l2_p0_col14_sum;
	
	assign comp_l2_p0_col15_cout = u_comp_l2_p0_col15_cout;
	
	assign comp_l2_p0_col15_sum = u_comp_l2_p0_col15_sum;
	
	assign comp_l2_p0_col16_cout = u_comp_l2_p0_col16_cout;
	
	assign comp_l2_p0_col16_sum = u_comp_l2_p0_col16_sum;
	
	assign comp_l2_p0_col17_cout = u_comp_l2_p0_col17_cout;
	
	assign comp_l2_p0_col17_sum = u_comp_l2_p0_col17_sum;
	
	assign comp_l2_p0_col18_cout = u_comp_l2_p0_col18_cout;
	
	assign comp_l2_p0_col18_sum = u_comp_l2_p0_col18_sum;
	
	assign comp_l2_p0_col19_cout = u_comp_l2_p0_col19_cout;
	
	assign comp_l2_p0_col19_sum = u_comp_l2_p0_col19_sum;
	
	assign comp_l2_p0_col20_cout = u_comp_l2_p0_col20_cout;
	
	assign comp_l2_p0_col20_sum = u_comp_l2_p0_col20_sum;
	
	assign comp_l2_p0_col21_cout = u_comp_l2_p0_col21_cout;
	
	assign comp_l2_p0_col21_sum = u_comp_l2_p0_col21_sum;
	
	assign comp_l2_p0_col22_cout = u_comp_l2_p0_col22_cout;
	
	assign comp_l2_p0_col22_sum = u_comp_l2_p0_col22_sum;
	
	assign comp_l2_p0_col23_cout = u_comp_l2_p0_col23_cout;
	
	assign comp_l2_p0_col23_sum = u_comp_l2_p0_col23_sum;
	
	assign comp_l2_p0_col24_cout = u_comp_l2_p0_col24_cout;
	
	assign comp_l2_p0_col24_sum = u_comp_l2_p0_col24_sum;
	
	assign comp_l2_p0_col25_cout = u_comp_l2_p0_col25_cout;
	
	assign comp_l2_p0_col25_sum = u_comp_l2_p0_col25_sum;
	
	assign comp_l2_p0_col26_cout = u_comp_l2_p0_col26_cout;
	
	assign comp_l2_p0_col26_sum = u_comp_l2_p0_col26_sum;
	
	assign comp_l2_p0_col27_cout = u_comp_l2_p0_col27_cout;
	
	assign comp_l2_p0_col27_sum = u_comp_l2_p0_col27_sum;
	
	assign comp_l2_p0_col28_cout = u_comp_l2_p0_col28_cout;
	
	assign comp_l2_p0_col28_sum = u_comp_l2_p0_col28_sum;
	
	assign comp_l2_p0_col29_cout = u_comp_l2_p0_col29_cout;
	
	assign comp_l2_p0_col29_sum = u_comp_l2_p0_col29_sum;
	
	assign comp_l2_p0_col30_cout = u_comp_l2_p0_col30_cout;
	
	assign comp_l2_p0_col30_sum = u_comp_l2_p0_col30_sum;
	
	assign comp_l2_p0_col31_sum = u_comp_l2_p0_col31_sum;
	
	assign comp_pad_l2_p0 = 1'b0;
	
	assign comp_l3_p0_col0_cout = u_comp_l3_p0_col0_cout;
	
	assign comp_l3_p0_col0_sum = u_comp_l3_p0_col0_sum;
	
	assign comp_l3_p0_col1_cout = u_comp_l3_p0_col1_cout;
	
	assign comp_l3_p0_col1_sum = u_comp_l3_p0_col1_sum;
	
	assign comp_l3_p0_col2_cout = u_comp_l3_p0_col2_cout;
	
	assign comp_l3_p0_col2_sum = u_comp_l3_p0_col2_sum;
	
	assign comp_l3_p0_col3_cout = u_comp_l3_p0_col3_cout;
	
	assign comp_l3_p0_col3_sum = u_comp_l3_p0_col3_sum;
	
	assign comp_l3_p0_col4_cout = u_comp_l3_p0_col4_cout;
	
	assign comp_l3_p0_col4_sum = u_comp_l3_p0_col4_sum;
	
	assign comp_l3_p0_col5_cout = u_comp_l3_p0_col5_cout;
	
	assign comp_l3_p0_col5_sum = u_comp_l3_p0_col5_sum;
	
	assign comp_l3_p0_col6_cout = u_comp_l3_p0_col6_cout;
	
	assign comp_l3_p0_col6_sum = u_comp_l3_p0_col6_sum;
	
	assign comp_l3_p0_col7_cout = u_comp_l3_p0_col7_cout;
	
	assign comp_l3_p0_col7_sum = u_comp_l3_p0_col7_sum;
	
	assign comp_l3_p0_col8_cout = u_comp_l3_p0_col8_cout;
	
	assign comp_l3_p0_col8_sum = u_comp_l3_p0_col8_sum;
	
	assign comp_l3_p0_col9_cout = u_comp_l3_p0_col9_cout;
	
	assign comp_l3_p0_col9_sum = u_comp_l3_p0_col9_sum;
	
	assign comp_l3_p0_col10_cout = u_comp_l3_p0_col10_cout;
	
	assign comp_l3_p0_col10_sum = u_comp_l3_p0_col10_sum;
	
	assign comp_l3_p0_col11_cout = u_comp_l3_p0_col11_cout;
	
	assign comp_l3_p0_col11_sum = u_comp_l3_p0_col11_sum;
	
	assign comp_l3_p0_col12_cout = u_comp_l3_p0_col12_cout;
	
	assign comp_l3_p0_col12_sum = u_comp_l3_p0_col12_sum;
	
	assign comp_l3_p0_col13_cout = u_comp_l3_p0_col13_cout;
	
	assign comp_l3_p0_col13_sum = u_comp_l3_p0_col13_sum;
	
	assign comp_l3_p0_col14_cout = u_comp_l3_p0_col14_cout;
	
	assign comp_l3_p0_col14_sum = u_comp_l3_p0_col14_sum;
	
	assign comp_l3_p0_col15_cout = u_comp_l3_p0_col15_cout;
	
	assign comp_l3_p0_col15_sum = u_comp_l3_p0_col15_sum;
	
	assign comp_l3_p0_col16_cout = u_comp_l3_p0_col16_cout;
	
	assign comp_l3_p0_col16_sum = u_comp_l3_p0_col16_sum;
	
	assign comp_l3_p0_col17_cout = u_comp_l3_p0_col17_cout;
	
	assign comp_l3_p0_col17_sum = u_comp_l3_p0_col17_sum;
	
	assign comp_l3_p0_col18_cout = u_comp_l3_p0_col18_cout;
	
	assign comp_l3_p0_col18_sum = u_comp_l3_p0_col18_sum;
	
	assign comp_l3_p0_col19_cout = u_comp_l3_p0_col19_cout;
	
	assign comp_l3_p0_col19_sum = u_comp_l3_p0_col19_sum;
	
	assign comp_l3_p0_col20_cout = u_comp_l3_p0_col20_cout;
	
	assign comp_l3_p0_col20_sum = u_comp_l3_p0_col20_sum;
	
	assign comp_l3_p0_col21_cout = u_comp_l3_p0_col21_cout;
	
	assign comp_l3_p0_col21_sum = u_comp_l3_p0_col21_sum;
	
	assign comp_l3_p0_col22_cout = u_comp_l3_p0_col22_cout;
	
	assign comp_l3_p0_col22_sum = u_comp_l3_p0_col22_sum;
	
	assign comp_l3_p0_col23_cout = u_comp_l3_p0_col23_cout;
	
	assign comp_l3_p0_col23_sum = u_comp_l3_p0_col23_sum;
	
	assign comp_l3_p0_col24_cout = u_comp_l3_p0_col24_cout;
	
	assign comp_l3_p0_col24_sum = u_comp_l3_p0_col24_sum;
	
	assign comp_l3_p0_col25_cout = u_comp_l3_p0_col25_cout;
	
	assign comp_l3_p0_col25_sum = u_comp_l3_p0_col25_sum;
	
	assign comp_l3_p0_col26_cout = u_comp_l3_p0_col26_cout;
	
	assign comp_l3_p0_col26_sum = u_comp_l3_p0_col26_sum;
	
	assign comp_l3_p0_col27_cout = u_comp_l3_p0_col27_cout;
	
	assign comp_l3_p0_col27_sum = u_comp_l3_p0_col27_sum;
	
	assign comp_l3_p0_col28_cout = u_comp_l3_p0_col28_cout;
	
	assign comp_l3_p0_col28_sum = u_comp_l3_p0_col28_sum;
	
	assign comp_l3_p0_col29_cout = u_comp_l3_p0_col29_cout;
	
	assign comp_l3_p0_col29_sum = u_comp_l3_p0_col29_sum;
	
	assign comp_l3_p0_col30_cout = u_comp_l3_p0_col30_cout;
	
	assign comp_l3_p0_col30_sum = u_comp_l3_p0_col30_sum;
	
	assign comp_l3_p0_col31_sum = u_comp_l3_p0_col31_sum;
	
	assign comp_pad_l3_p0 = 1'b0;
	
	assign comp_l4_p0_col0_cout = u_comp_l4_p0_col0_cout;
	
	assign comp_l4_p0_col0_sum = u_comp_l4_p0_col0_sum;
	
	assign comp_l4_p0_col1_cout = u_comp_l4_p0_col1_cout;
	
	assign comp_l4_p0_col1_sum = u_comp_l4_p0_col1_sum;
	
	assign comp_l4_p0_col2_cout = u_comp_l4_p0_col2_cout;
	
	assign comp_l4_p0_col2_sum = u_comp_l4_p0_col2_sum;
	
	assign comp_l4_p0_col3_cout = u_comp_l4_p0_col3_cout;
	
	assign comp_l4_p0_col3_sum = u_comp_l4_p0_col3_sum;
	
	assign comp_l4_p0_col4_cout = u_comp_l4_p0_col4_cout;
	
	assign comp_l4_p0_col4_sum = u_comp_l4_p0_col4_sum;
	
	assign comp_l4_p0_col5_cout = u_comp_l4_p0_col5_cout;
	
	assign comp_l4_p0_col5_sum = u_comp_l4_p0_col5_sum;
	
	assign comp_l4_p0_col6_cout = u_comp_l4_p0_col6_cout;
	
	assign comp_l4_p0_col6_sum = u_comp_l4_p0_col6_sum;
	
	assign comp_l4_p0_col7_cout = u_comp_l4_p0_col7_cout;
	
	assign comp_l4_p0_col7_sum = u_comp_l4_p0_col7_sum;
	
	assign comp_l4_p0_col8_cout = u_comp_l4_p0_col8_cout;
	
	assign comp_l4_p0_col8_sum = u_comp_l4_p0_col8_sum;
	
	assign comp_l4_p0_col9_cout = u_comp_l4_p0_col9_cout;
	
	assign comp_l4_p0_col9_sum = u_comp_l4_p0_col9_sum;
	
	assign comp_l4_p0_col10_cout = u_comp_l4_p0_col10_cout;
	
	assign comp_l4_p0_col10_sum = u_comp_l4_p0_col10_sum;
	
	assign comp_l4_p0_col11_cout = u_comp_l4_p0_col11_cout;
	
	assign comp_l4_p0_col11_sum = u_comp_l4_p0_col11_sum;
	
	assign comp_l4_p0_col12_cout = u_comp_l4_p0_col12_cout;
	
	assign comp_l4_p0_col12_sum = u_comp_l4_p0_col12_sum;
	
	assign comp_l4_p0_col13_cout = u_comp_l4_p0_col13_cout;
	
	assign comp_l4_p0_col13_sum = u_comp_l4_p0_col13_sum;
	
	assign comp_l4_p0_col14_cout = u_comp_l4_p0_col14_cout;
	
	assign comp_l4_p0_col14_sum = u_comp_l4_p0_col14_sum;
	
	assign comp_l4_p0_col15_cout = u_comp_l4_p0_col15_cout;
	
	assign comp_l4_p0_col15_sum = u_comp_l4_p0_col15_sum;
	
	assign comp_l4_p0_col16_cout = u_comp_l4_p0_col16_cout;
	
	assign comp_l4_p0_col16_sum = u_comp_l4_p0_col16_sum;
	
	assign comp_l4_p0_col17_cout = u_comp_l4_p0_col17_cout;
	
	assign comp_l4_p0_col17_sum = u_comp_l4_p0_col17_sum;
	
	assign comp_l4_p0_col18_cout = u_comp_l4_p0_col18_cout;
	
	assign comp_l4_p0_col18_sum = u_comp_l4_p0_col18_sum;
	
	assign comp_l4_p0_col19_cout = u_comp_l4_p0_col19_cout;
	
	assign comp_l4_p0_col19_sum = u_comp_l4_p0_col19_sum;
	
	assign comp_l4_p0_col20_cout = u_comp_l4_p0_col20_cout;
	
	assign comp_l4_p0_col20_sum = u_comp_l4_p0_col20_sum;
	
	assign comp_l4_p0_col21_cout = u_comp_l4_p0_col21_cout;
	
	assign comp_l4_p0_col21_sum = u_comp_l4_p0_col21_sum;
	
	assign comp_l4_p0_col22_cout = u_comp_l4_p0_col22_cout;
	
	assign comp_l4_p0_col22_sum = u_comp_l4_p0_col22_sum;
	
	assign comp_l4_p0_col23_cout = u_comp_l4_p0_col23_cout;
	
	assign comp_l4_p0_col23_sum = u_comp_l4_p0_col23_sum;
	
	assign comp_l4_p0_col24_cout = u_comp_l4_p0_col24_cout;
	
	assign comp_l4_p0_col24_sum = u_comp_l4_p0_col24_sum;
	
	assign comp_l4_p0_col25_cout = u_comp_l4_p0_col25_cout;
	
	assign comp_l4_p0_col25_sum = u_comp_l4_p0_col25_sum;
	
	assign comp_l4_p0_col26_cout = u_comp_l4_p0_col26_cout;
	
	assign comp_l4_p0_col26_sum = u_comp_l4_p0_col26_sum;
	
	assign comp_l4_p0_col27_cout = u_comp_l4_p0_col27_cout;
	
	assign comp_l4_p0_col27_sum = u_comp_l4_p0_col27_sum;
	
	assign comp_l4_p0_col28_cout = u_comp_l4_p0_col28_cout;
	
	assign comp_l4_p0_col28_sum = u_comp_l4_p0_col28_sum;
	
	assign comp_l4_p0_col29_cout = u_comp_l4_p0_col29_cout;
	
	assign comp_l4_p0_col29_sum = u_comp_l4_p0_col29_sum;
	
	assign comp_l4_p0_col30_cout = u_comp_l4_p0_col30_cout;
	
	assign comp_l4_p0_col30_sum = u_comp_l4_p0_col30_sum;
	
	assign comp_l4_p0_col31_sum = u_comp_l4_p0_col31_sum;
	
	assign comp_pad_l4_p0 = 1'b0;
	

	//Wire this module connect to sub module.
	assign u_comp_l0_p0_col0_a = p_0_0;
	
	assign u_comp_l0_p0_col0_b = p_1_0;
	
	assign u_comp_l0_p0_col0_cin = p_2_0;
	
	assign u_comp_l0_p0_col1_a = p_0_1;
	
	assign u_comp_l0_p0_col1_b = p_1_1;
	
	assign u_comp_l0_p0_col1_cin = p_2_1;
	
	assign u_comp_l0_p0_col2_a = p_0_2;
	
	assign u_comp_l0_p0_col2_b = p_1_2;
	
	assign u_comp_l0_p0_col2_cin = p_2_2;
	
	assign u_comp_l0_p0_col3_a = p_0_3;
	
	assign u_comp_l0_p0_col3_b = p_1_3;
	
	assign u_comp_l0_p0_col3_cin = p_2_3;
	
	assign u_comp_l0_p0_col4_a = p_0_4;
	
	assign u_comp_l0_p0_col4_b = p_1_4;
	
	assign u_comp_l0_p0_col4_cin = p_2_4;
	
	assign u_comp_l0_p0_col5_a = p_0_5;
	
	assign u_comp_l0_p0_col5_b = p_1_5;
	
	assign u_comp_l0_p0_col5_cin = p_2_5;
	
	assign u_comp_l0_p0_col6_a = p_0_6;
	
	assign u_comp_l0_p0_col6_b = p_1_6;
	
	assign u_comp_l0_p0_col6_cin = p_2_6;
	
	assign u_comp_l0_p0_col7_a = p_0_7;
	
	assign u_comp_l0_p0_col7_b = p_1_7;
	
	assign u_comp_l0_p0_col7_cin = p_2_7;
	
	assign u_comp_l0_p0_col8_a = p_0_8;
	
	assign u_comp_l0_p0_col8_b = p_1_8;
	
	assign u_comp_l0_p0_col8_cin = p_2_8;
	
	assign u_comp_l0_p0_col9_a = p_0_9;
	
	assign u_comp_l0_p0_col9_b = p_1_9;
	
	assign u_comp_l0_p0_col9_cin = p_2_9;
	
	assign u_comp_l0_p0_col10_a = p_0_10;
	
	assign u_comp_l0_p0_col10_b = p_1_10;
	
	assign u_comp_l0_p0_col10_cin = p_2_10;
	
	assign u_comp_l0_p0_col11_a = p_0_11;
	
	assign u_comp_l0_p0_col11_b = p_1_11;
	
	assign u_comp_l0_p0_col11_cin = p_2_11;
	
	assign u_comp_l0_p0_col12_a = p_0_12;
	
	assign u_comp_l0_p0_col12_b = p_1_12;
	
	assign u_comp_l0_p0_col12_cin = p_2_12;
	
	assign u_comp_l0_p0_col13_a = p_0_13;
	
	assign u_comp_l0_p0_col13_b = p_1_13;
	
	assign u_comp_l0_p0_col13_cin = p_2_13;
	
	assign u_comp_l0_p0_col14_a = p_0_14;
	
	assign u_comp_l0_p0_col14_b = p_1_14;
	
	assign u_comp_l0_p0_col14_cin = p_2_14;
	
	assign u_comp_l0_p0_col15_a = p_0_15;
	
	assign u_comp_l0_p0_col15_b = p_1_15;
	
	assign u_comp_l0_p0_col15_cin = p_2_15;
	
	assign u_comp_l0_p0_col16_a = p_0_16;
	
	assign u_comp_l0_p0_col16_b = p_1_16;
	
	assign u_comp_l0_p0_col16_cin = p_2_16;
	
	assign u_comp_l0_p0_col17_a = p_0_17;
	
	assign u_comp_l0_p0_col17_b = p_1_17;
	
	assign u_comp_l0_p0_col17_cin = p_2_17;
	
	assign u_comp_l0_p0_col18_a = p_0_18;
	
	assign u_comp_l0_p0_col18_b = p_1_18;
	
	assign u_comp_l0_p0_col18_cin = p_2_18;
	
	assign u_comp_l0_p0_col19_a = p_0_19;
	
	assign u_comp_l0_p0_col19_b = p_1_19;
	
	assign u_comp_l0_p0_col19_cin = p_2_19;
	
	assign u_comp_l0_p0_col20_a = p_0_20;
	
	assign u_comp_l0_p0_col20_b = p_1_20;
	
	assign u_comp_l0_p0_col20_cin = p_2_20;
	
	assign u_comp_l0_p0_col21_a = p_0_21;
	
	assign u_comp_l0_p0_col21_b = p_1_21;
	
	assign u_comp_l0_p0_col21_cin = p_2_21;
	
	assign u_comp_l0_p0_col22_a = p_0_22;
	
	assign u_comp_l0_p0_col22_b = p_1_22;
	
	assign u_comp_l0_p0_col22_cin = p_2_22;
	
	assign u_comp_l0_p0_col23_a = p_0_23;
	
	assign u_comp_l0_p0_col23_b = p_1_23;
	
	assign u_comp_l0_p0_col23_cin = p_2_23;
	
	assign u_comp_l0_p0_col24_a = p_0_24;
	
	assign u_comp_l0_p0_col24_b = p_1_24;
	
	assign u_comp_l0_p0_col24_cin = p_2_24;
	
	assign u_comp_l0_p0_col25_a = p_0_25;
	
	assign u_comp_l0_p0_col25_b = p_1_25;
	
	assign u_comp_l0_p0_col25_cin = p_2_25;
	
	assign u_comp_l0_p0_col26_a = p_0_26;
	
	assign u_comp_l0_p0_col26_b = p_1_26;
	
	assign u_comp_l0_p0_col26_cin = p_2_26;
	
	assign u_comp_l0_p0_col27_a = p_0_27;
	
	assign u_comp_l0_p0_col27_b = p_1_27;
	
	assign u_comp_l0_p0_col27_cin = p_2_27;
	
	assign u_comp_l0_p0_col28_a = p_0_28;
	
	assign u_comp_l0_p0_col28_b = p_1_28;
	
	assign u_comp_l0_p0_col28_cin = p_2_28;
	
	assign u_comp_l0_p0_col29_a = p_0_29;
	
	assign u_comp_l0_p0_col29_b = p_1_29;
	
	assign u_comp_l0_p0_col29_cin = p_2_29;
	
	assign u_comp_l0_p0_col30_a = p_0_30;
	
	assign u_comp_l0_p0_col30_b = p_1_30;
	
	assign u_comp_l0_p0_col30_cin = p_2_30;
	
	assign u_comp_l0_p0_col31_a = p_0_31;
	
	assign u_comp_l0_p0_col31_b = p_1_31;
	
	assign u_comp_l0_p0_col31_cin = p_2_31;
	
	assign u_comp_l0_p1_col0_a = p_3_0;
	
	assign u_comp_l0_p1_col0_b = p_4_0;
	
	assign u_comp_l0_p1_col0_cin = p_5_0;
	
	assign u_comp_l0_p1_col1_a = p_3_1;
	
	assign u_comp_l0_p1_col1_b = p_4_1;
	
	assign u_comp_l0_p1_col1_cin = p_5_1;
	
	assign u_comp_l0_p1_col2_a = p_3_2;
	
	assign u_comp_l0_p1_col2_b = p_4_2;
	
	assign u_comp_l0_p1_col2_cin = p_5_2;
	
	assign u_comp_l0_p1_col3_a = p_3_3;
	
	assign u_comp_l0_p1_col3_b = p_4_3;
	
	assign u_comp_l0_p1_col3_cin = p_5_3;
	
	assign u_comp_l0_p1_col4_a = p_3_4;
	
	assign u_comp_l0_p1_col4_b = p_4_4;
	
	assign u_comp_l0_p1_col4_cin = p_5_4;
	
	assign u_comp_l0_p1_col5_a = p_3_5;
	
	assign u_comp_l0_p1_col5_b = p_4_5;
	
	assign u_comp_l0_p1_col5_cin = p_5_5;
	
	assign u_comp_l0_p1_col6_a = p_3_6;
	
	assign u_comp_l0_p1_col6_b = p_4_6;
	
	assign u_comp_l0_p1_col6_cin = p_5_6;
	
	assign u_comp_l0_p1_col7_a = p_3_7;
	
	assign u_comp_l0_p1_col7_b = p_4_7;
	
	assign u_comp_l0_p1_col7_cin = p_5_7;
	
	assign u_comp_l0_p1_col8_a = p_3_8;
	
	assign u_comp_l0_p1_col8_b = p_4_8;
	
	assign u_comp_l0_p1_col8_cin = p_5_8;
	
	assign u_comp_l0_p1_col9_a = p_3_9;
	
	assign u_comp_l0_p1_col9_b = p_4_9;
	
	assign u_comp_l0_p1_col9_cin = p_5_9;
	
	assign u_comp_l0_p1_col10_a = p_3_10;
	
	assign u_comp_l0_p1_col10_b = p_4_10;
	
	assign u_comp_l0_p1_col10_cin = p_5_10;
	
	assign u_comp_l0_p1_col11_a = p_3_11;
	
	assign u_comp_l0_p1_col11_b = p_4_11;
	
	assign u_comp_l0_p1_col11_cin = p_5_11;
	
	assign u_comp_l0_p1_col12_a = p_3_12;
	
	assign u_comp_l0_p1_col12_b = p_4_12;
	
	assign u_comp_l0_p1_col12_cin = p_5_12;
	
	assign u_comp_l0_p1_col13_a = p_3_13;
	
	assign u_comp_l0_p1_col13_b = p_4_13;
	
	assign u_comp_l0_p1_col13_cin = p_5_13;
	
	assign u_comp_l0_p1_col14_a = p_3_14;
	
	assign u_comp_l0_p1_col14_b = p_4_14;
	
	assign u_comp_l0_p1_col14_cin = p_5_14;
	
	assign u_comp_l0_p1_col15_a = p_3_15;
	
	assign u_comp_l0_p1_col15_b = p_4_15;
	
	assign u_comp_l0_p1_col15_cin = p_5_15;
	
	assign u_comp_l0_p1_col16_a = p_3_16;
	
	assign u_comp_l0_p1_col16_b = p_4_16;
	
	assign u_comp_l0_p1_col16_cin = p_5_16;
	
	assign u_comp_l0_p1_col17_a = p_3_17;
	
	assign u_comp_l0_p1_col17_b = p_4_17;
	
	assign u_comp_l0_p1_col17_cin = p_5_17;
	
	assign u_comp_l0_p1_col18_a = p_3_18;
	
	assign u_comp_l0_p1_col18_b = p_4_18;
	
	assign u_comp_l0_p1_col18_cin = p_5_18;
	
	assign u_comp_l0_p1_col19_a = p_3_19;
	
	assign u_comp_l0_p1_col19_b = p_4_19;
	
	assign u_comp_l0_p1_col19_cin = p_5_19;
	
	assign u_comp_l0_p1_col20_a = p_3_20;
	
	assign u_comp_l0_p1_col20_b = p_4_20;
	
	assign u_comp_l0_p1_col20_cin = p_5_20;
	
	assign u_comp_l0_p1_col21_a = p_3_21;
	
	assign u_comp_l0_p1_col21_b = p_4_21;
	
	assign u_comp_l0_p1_col21_cin = p_5_21;
	
	assign u_comp_l0_p1_col22_a = p_3_22;
	
	assign u_comp_l0_p1_col22_b = p_4_22;
	
	assign u_comp_l0_p1_col22_cin = p_5_22;
	
	assign u_comp_l0_p1_col23_a = p_3_23;
	
	assign u_comp_l0_p1_col23_b = p_4_23;
	
	assign u_comp_l0_p1_col23_cin = p_5_23;
	
	assign u_comp_l0_p1_col24_a = p_3_24;
	
	assign u_comp_l0_p1_col24_b = p_4_24;
	
	assign u_comp_l0_p1_col24_cin = p_5_24;
	
	assign u_comp_l0_p1_col25_a = p_3_25;
	
	assign u_comp_l0_p1_col25_b = p_4_25;
	
	assign u_comp_l0_p1_col25_cin = p_5_25;
	
	assign u_comp_l0_p1_col26_a = p_3_26;
	
	assign u_comp_l0_p1_col26_b = p_4_26;
	
	assign u_comp_l0_p1_col26_cin = p_5_26;
	
	assign u_comp_l0_p1_col27_a = p_3_27;
	
	assign u_comp_l0_p1_col27_b = p_4_27;
	
	assign u_comp_l0_p1_col27_cin = p_5_27;
	
	assign u_comp_l0_p1_col28_a = p_3_28;
	
	assign u_comp_l0_p1_col28_b = p_4_28;
	
	assign u_comp_l0_p1_col28_cin = p_5_28;
	
	assign u_comp_l0_p1_col29_a = p_3_29;
	
	assign u_comp_l0_p1_col29_b = p_4_29;
	
	assign u_comp_l0_p1_col29_cin = p_5_29;
	
	assign u_comp_l0_p1_col30_a = p_3_30;
	
	assign u_comp_l0_p1_col30_b = p_4_30;
	
	assign u_comp_l0_p1_col30_cin = p_5_30;
	
	assign u_comp_l0_p1_col31_a = p_3_31;
	
	assign u_comp_l0_p1_col31_b = p_4_31;
	
	assign u_comp_l0_p1_col31_cin = p_5_31;
	
	assign u_comp_l0_p2_col0_a = p_6_0;
	
	assign u_comp_l0_p2_col0_b = p_7_0;
	
	assign u_comp_l0_p2_col0_cin = p_8_0;
	
	assign u_comp_l0_p2_col1_a = p_6_1;
	
	assign u_comp_l0_p2_col1_b = p_7_1;
	
	assign u_comp_l0_p2_col1_cin = p_8_1;
	
	assign u_comp_l0_p2_col2_a = p_6_2;
	
	assign u_comp_l0_p2_col2_b = p_7_2;
	
	assign u_comp_l0_p2_col2_cin = p_8_2;
	
	assign u_comp_l0_p2_col3_a = p_6_3;
	
	assign u_comp_l0_p2_col3_b = p_7_3;
	
	assign u_comp_l0_p2_col3_cin = p_8_3;
	
	assign u_comp_l0_p2_col4_a = p_6_4;
	
	assign u_comp_l0_p2_col4_b = p_7_4;
	
	assign u_comp_l0_p2_col4_cin = p_8_4;
	
	assign u_comp_l0_p2_col5_a = p_6_5;
	
	assign u_comp_l0_p2_col5_b = p_7_5;
	
	assign u_comp_l0_p2_col5_cin = p_8_5;
	
	assign u_comp_l0_p2_col6_a = p_6_6;
	
	assign u_comp_l0_p2_col6_b = p_7_6;
	
	assign u_comp_l0_p2_col6_cin = p_8_6;
	
	assign u_comp_l0_p2_col7_a = p_6_7;
	
	assign u_comp_l0_p2_col7_b = p_7_7;
	
	assign u_comp_l0_p2_col7_cin = p_8_7;
	
	assign u_comp_l0_p2_col8_a = p_6_8;
	
	assign u_comp_l0_p2_col8_b = p_7_8;
	
	assign u_comp_l0_p2_col8_cin = p_8_8;
	
	assign u_comp_l0_p2_col9_a = p_6_9;
	
	assign u_comp_l0_p2_col9_b = p_7_9;
	
	assign u_comp_l0_p2_col9_cin = p_8_9;
	
	assign u_comp_l0_p2_col10_a = p_6_10;
	
	assign u_comp_l0_p2_col10_b = p_7_10;
	
	assign u_comp_l0_p2_col10_cin = p_8_10;
	
	assign u_comp_l0_p2_col11_a = p_6_11;
	
	assign u_comp_l0_p2_col11_b = p_7_11;
	
	assign u_comp_l0_p2_col11_cin = p_8_11;
	
	assign u_comp_l0_p2_col12_a = p_6_12;
	
	assign u_comp_l0_p2_col12_b = p_7_12;
	
	assign u_comp_l0_p2_col12_cin = p_8_12;
	
	assign u_comp_l0_p2_col13_a = p_6_13;
	
	assign u_comp_l0_p2_col13_b = p_7_13;
	
	assign u_comp_l0_p2_col13_cin = p_8_13;
	
	assign u_comp_l0_p2_col14_a = p_6_14;
	
	assign u_comp_l0_p2_col14_b = p_7_14;
	
	assign u_comp_l0_p2_col14_cin = p_8_14;
	
	assign u_comp_l0_p2_col15_a = p_6_15;
	
	assign u_comp_l0_p2_col15_b = p_7_15;
	
	assign u_comp_l0_p2_col15_cin = p_8_15;
	
	assign u_comp_l0_p2_col16_a = p_6_16;
	
	assign u_comp_l0_p2_col16_b = p_7_16;
	
	assign u_comp_l0_p2_col16_cin = p_8_16;
	
	assign u_comp_l0_p2_col17_a = p_6_17;
	
	assign u_comp_l0_p2_col17_b = p_7_17;
	
	assign u_comp_l0_p2_col17_cin = p_8_17;
	
	assign u_comp_l0_p2_col18_a = p_6_18;
	
	assign u_comp_l0_p2_col18_b = p_7_18;
	
	assign u_comp_l0_p2_col18_cin = p_8_18;
	
	assign u_comp_l0_p2_col19_a = p_6_19;
	
	assign u_comp_l0_p2_col19_b = p_7_19;
	
	assign u_comp_l0_p2_col19_cin = p_8_19;
	
	assign u_comp_l0_p2_col20_a = p_6_20;
	
	assign u_comp_l0_p2_col20_b = p_7_20;
	
	assign u_comp_l0_p2_col20_cin = p_8_20;
	
	assign u_comp_l0_p2_col21_a = p_6_21;
	
	assign u_comp_l0_p2_col21_b = p_7_21;
	
	assign u_comp_l0_p2_col21_cin = p_8_21;
	
	assign u_comp_l0_p2_col22_a = p_6_22;
	
	assign u_comp_l0_p2_col22_b = p_7_22;
	
	assign u_comp_l0_p2_col22_cin = p_8_22;
	
	assign u_comp_l0_p2_col23_a = p_6_23;
	
	assign u_comp_l0_p2_col23_b = p_7_23;
	
	assign u_comp_l0_p2_col23_cin = p_8_23;
	
	assign u_comp_l0_p2_col24_a = p_6_24;
	
	assign u_comp_l0_p2_col24_b = p_7_24;
	
	assign u_comp_l0_p2_col24_cin = p_8_24;
	
	assign u_comp_l0_p2_col25_a = p_6_25;
	
	assign u_comp_l0_p2_col25_b = p_7_25;
	
	assign u_comp_l0_p2_col25_cin = p_8_25;
	
	assign u_comp_l0_p2_col26_a = p_6_26;
	
	assign u_comp_l0_p2_col26_b = p_7_26;
	
	assign u_comp_l0_p2_col26_cin = p_8_26;
	
	assign u_comp_l0_p2_col27_a = p_6_27;
	
	assign u_comp_l0_p2_col27_b = p_7_27;
	
	assign u_comp_l0_p2_col27_cin = p_8_27;
	
	assign u_comp_l0_p2_col28_a = p_6_28;
	
	assign u_comp_l0_p2_col28_b = p_7_28;
	
	assign u_comp_l0_p2_col28_cin = p_8_28;
	
	assign u_comp_l0_p2_col29_a = p_6_29;
	
	assign u_comp_l0_p2_col29_b = p_7_29;
	
	assign u_comp_l0_p2_col29_cin = p_8_29;
	
	assign u_comp_l0_p2_col30_a = p_6_30;
	
	assign u_comp_l0_p2_col30_b = p_7_30;
	
	assign u_comp_l0_p2_col30_cin = p_8_30;
	
	assign u_comp_l0_p2_col31_a = p_6_31;
	
	assign u_comp_l0_p2_col31_b = p_7_31;
	
	assign u_comp_l0_p2_col31_cin = p_8_31;
	
	assign u_comp_l1_p0_col0_a = comp_l0_p0_col0_sum;
	
	assign u_comp_l1_p0_col0_b = comp_pad_l0_p0;
	
	assign u_comp_l1_p0_col0_cin = comp_l0_p1_col0_sum;
	
	assign u_comp_l1_p0_col1_a = comp_l0_p0_col1_sum;
	
	assign u_comp_l1_p0_col1_b = comp_l0_p0_col0_cout;
	
	assign u_comp_l1_p0_col1_cin = comp_l0_p1_col1_sum;
	
	assign u_comp_l1_p0_col2_a = comp_l0_p0_col2_sum;
	
	assign u_comp_l1_p0_col2_b = comp_l0_p0_col1_cout;
	
	assign u_comp_l1_p0_col2_cin = comp_l0_p1_col2_sum;
	
	assign u_comp_l1_p0_col3_a = comp_l0_p0_col3_sum;
	
	assign u_comp_l1_p0_col3_b = comp_l0_p0_col2_cout;
	
	assign u_comp_l1_p0_col3_cin = comp_l0_p1_col3_sum;
	
	assign u_comp_l1_p0_col4_a = comp_l0_p0_col4_sum;
	
	assign u_comp_l1_p0_col4_b = comp_l0_p0_col3_cout;
	
	assign u_comp_l1_p0_col4_cin = comp_l0_p1_col4_sum;
	
	assign u_comp_l1_p0_col5_a = comp_l0_p0_col5_sum;
	
	assign u_comp_l1_p0_col5_b = comp_l0_p0_col4_cout;
	
	assign u_comp_l1_p0_col5_cin = comp_l0_p1_col5_sum;
	
	assign u_comp_l1_p0_col6_a = comp_l0_p0_col6_sum;
	
	assign u_comp_l1_p0_col6_b = comp_l0_p0_col5_cout;
	
	assign u_comp_l1_p0_col6_cin = comp_l0_p1_col6_sum;
	
	assign u_comp_l1_p0_col7_a = comp_l0_p0_col7_sum;
	
	assign u_comp_l1_p0_col7_b = comp_l0_p0_col6_cout;
	
	assign u_comp_l1_p0_col7_cin = comp_l0_p1_col7_sum;
	
	assign u_comp_l1_p0_col8_a = comp_l0_p0_col8_sum;
	
	assign u_comp_l1_p0_col8_b = comp_l0_p0_col7_cout;
	
	assign u_comp_l1_p0_col8_cin = comp_l0_p1_col8_sum;
	
	assign u_comp_l1_p0_col9_a = comp_l0_p0_col9_sum;
	
	assign u_comp_l1_p0_col9_b = comp_l0_p0_col8_cout;
	
	assign u_comp_l1_p0_col9_cin = comp_l0_p1_col9_sum;
	
	assign u_comp_l1_p0_col10_a = comp_l0_p0_col10_sum;
	
	assign u_comp_l1_p0_col10_b = comp_l0_p0_col9_cout;
	
	assign u_comp_l1_p0_col10_cin = comp_l0_p1_col10_sum;
	
	assign u_comp_l1_p0_col11_a = comp_l0_p0_col11_sum;
	
	assign u_comp_l1_p0_col11_b = comp_l0_p0_col10_cout;
	
	assign u_comp_l1_p0_col11_cin = comp_l0_p1_col11_sum;
	
	assign u_comp_l1_p0_col12_a = comp_l0_p0_col12_sum;
	
	assign u_comp_l1_p0_col12_b = comp_l0_p0_col11_cout;
	
	assign u_comp_l1_p0_col12_cin = comp_l0_p1_col12_sum;
	
	assign u_comp_l1_p0_col13_a = comp_l0_p0_col13_sum;
	
	assign u_comp_l1_p0_col13_b = comp_l0_p0_col12_cout;
	
	assign u_comp_l1_p0_col13_cin = comp_l0_p1_col13_sum;
	
	assign u_comp_l1_p0_col14_a = comp_l0_p0_col14_sum;
	
	assign u_comp_l1_p0_col14_b = comp_l0_p0_col13_cout;
	
	assign u_comp_l1_p0_col14_cin = comp_l0_p1_col14_sum;
	
	assign u_comp_l1_p0_col15_a = comp_l0_p0_col15_sum;
	
	assign u_comp_l1_p0_col15_b = comp_l0_p0_col14_cout;
	
	assign u_comp_l1_p0_col15_cin = comp_l0_p1_col15_sum;
	
	assign u_comp_l1_p0_col16_a = comp_l0_p0_col16_sum;
	
	assign u_comp_l1_p0_col16_b = comp_l0_p0_col15_cout;
	
	assign u_comp_l1_p0_col16_cin = comp_l0_p1_col16_sum;
	
	assign u_comp_l1_p0_col17_a = comp_l0_p0_col17_sum;
	
	assign u_comp_l1_p0_col17_b = comp_l0_p0_col16_cout;
	
	assign u_comp_l1_p0_col17_cin = comp_l0_p1_col17_sum;
	
	assign u_comp_l1_p0_col18_a = comp_l0_p0_col18_sum;
	
	assign u_comp_l1_p0_col18_b = comp_l0_p0_col17_cout;
	
	assign u_comp_l1_p0_col18_cin = comp_l0_p1_col18_sum;
	
	assign u_comp_l1_p0_col19_a = comp_l0_p0_col19_sum;
	
	assign u_comp_l1_p0_col19_b = comp_l0_p0_col18_cout;
	
	assign u_comp_l1_p0_col19_cin = comp_l0_p1_col19_sum;
	
	assign u_comp_l1_p0_col20_a = comp_l0_p0_col20_sum;
	
	assign u_comp_l1_p0_col20_b = comp_l0_p0_col19_cout;
	
	assign u_comp_l1_p0_col20_cin = comp_l0_p1_col20_sum;
	
	assign u_comp_l1_p0_col21_a = comp_l0_p0_col21_sum;
	
	assign u_comp_l1_p0_col21_b = comp_l0_p0_col20_cout;
	
	assign u_comp_l1_p0_col21_cin = comp_l0_p1_col21_sum;
	
	assign u_comp_l1_p0_col22_a = comp_l0_p0_col22_sum;
	
	assign u_comp_l1_p0_col22_b = comp_l0_p0_col21_cout;
	
	assign u_comp_l1_p0_col22_cin = comp_l0_p1_col22_sum;
	
	assign u_comp_l1_p0_col23_a = comp_l0_p0_col23_sum;
	
	assign u_comp_l1_p0_col23_b = comp_l0_p0_col22_cout;
	
	assign u_comp_l1_p0_col23_cin = comp_l0_p1_col23_sum;
	
	assign u_comp_l1_p0_col24_a = comp_l0_p0_col24_sum;
	
	assign u_comp_l1_p0_col24_b = comp_l0_p0_col23_cout;
	
	assign u_comp_l1_p0_col24_cin = comp_l0_p1_col24_sum;
	
	assign u_comp_l1_p0_col25_a = comp_l0_p0_col25_sum;
	
	assign u_comp_l1_p0_col25_b = comp_l0_p0_col24_cout;
	
	assign u_comp_l1_p0_col25_cin = comp_l0_p1_col25_sum;
	
	assign u_comp_l1_p0_col26_a = comp_l0_p0_col26_sum;
	
	assign u_comp_l1_p0_col26_b = comp_l0_p0_col25_cout;
	
	assign u_comp_l1_p0_col26_cin = comp_l0_p1_col26_sum;
	
	assign u_comp_l1_p0_col27_a = comp_l0_p0_col27_sum;
	
	assign u_comp_l1_p0_col27_b = comp_l0_p0_col26_cout;
	
	assign u_comp_l1_p0_col27_cin = comp_l0_p1_col27_sum;
	
	assign u_comp_l1_p0_col28_a = comp_l0_p0_col28_sum;
	
	assign u_comp_l1_p0_col28_b = comp_l0_p0_col27_cout;
	
	assign u_comp_l1_p0_col28_cin = comp_l0_p1_col28_sum;
	
	assign u_comp_l1_p0_col29_a = comp_l0_p0_col29_sum;
	
	assign u_comp_l1_p0_col29_b = comp_l0_p0_col28_cout;
	
	assign u_comp_l1_p0_col29_cin = comp_l0_p1_col29_sum;
	
	assign u_comp_l1_p0_col30_a = comp_l0_p0_col30_sum;
	
	assign u_comp_l1_p0_col30_b = comp_l0_p0_col29_cout;
	
	assign u_comp_l1_p0_col30_cin = comp_l0_p1_col30_sum;
	
	assign u_comp_l1_p0_col31_a = comp_l0_p0_col31_sum;
	
	assign u_comp_l1_p0_col31_b = comp_l0_p0_col30_cout;
	
	assign u_comp_l1_p0_col31_cin = comp_l0_p1_col31_sum;
	
	assign u_comp_l1_p1_col0_a = comp_pad_l0_p1;
	
	assign u_comp_l1_p1_col0_b = comp_l0_p2_col0_sum;
	
	assign u_comp_l1_p1_col0_cin = comp_pad_l0_p2;
	
	assign u_comp_l1_p1_col1_a = comp_l0_p1_col0_cout;
	
	assign u_comp_l1_p1_col1_b = comp_l0_p2_col1_sum;
	
	assign u_comp_l1_p1_col1_cin = comp_l0_p2_col0_cout;
	
	assign u_comp_l1_p1_col2_a = comp_l0_p1_col1_cout;
	
	assign u_comp_l1_p1_col2_b = comp_l0_p2_col2_sum;
	
	assign u_comp_l1_p1_col2_cin = comp_l0_p2_col1_cout;
	
	assign u_comp_l1_p1_col3_a = comp_l0_p1_col2_cout;
	
	assign u_comp_l1_p1_col3_b = comp_l0_p2_col3_sum;
	
	assign u_comp_l1_p1_col3_cin = comp_l0_p2_col2_cout;
	
	assign u_comp_l1_p1_col4_a = comp_l0_p1_col3_cout;
	
	assign u_comp_l1_p1_col4_b = comp_l0_p2_col4_sum;
	
	assign u_comp_l1_p1_col4_cin = comp_l0_p2_col3_cout;
	
	assign u_comp_l1_p1_col5_a = comp_l0_p1_col4_cout;
	
	assign u_comp_l1_p1_col5_b = comp_l0_p2_col5_sum;
	
	assign u_comp_l1_p1_col5_cin = comp_l0_p2_col4_cout;
	
	assign u_comp_l1_p1_col6_a = comp_l0_p1_col5_cout;
	
	assign u_comp_l1_p1_col6_b = comp_l0_p2_col6_sum;
	
	assign u_comp_l1_p1_col6_cin = comp_l0_p2_col5_cout;
	
	assign u_comp_l1_p1_col7_a = comp_l0_p1_col6_cout;
	
	assign u_comp_l1_p1_col7_b = comp_l0_p2_col7_sum;
	
	assign u_comp_l1_p1_col7_cin = comp_l0_p2_col6_cout;
	
	assign u_comp_l1_p1_col8_a = comp_l0_p1_col7_cout;
	
	assign u_comp_l1_p1_col8_b = comp_l0_p2_col8_sum;
	
	assign u_comp_l1_p1_col8_cin = comp_l0_p2_col7_cout;
	
	assign u_comp_l1_p1_col9_a = comp_l0_p1_col8_cout;
	
	assign u_comp_l1_p1_col9_b = comp_l0_p2_col9_sum;
	
	assign u_comp_l1_p1_col9_cin = comp_l0_p2_col8_cout;
	
	assign u_comp_l1_p1_col10_a = comp_l0_p1_col9_cout;
	
	assign u_comp_l1_p1_col10_b = comp_l0_p2_col10_sum;
	
	assign u_comp_l1_p1_col10_cin = comp_l0_p2_col9_cout;
	
	assign u_comp_l1_p1_col11_a = comp_l0_p1_col10_cout;
	
	assign u_comp_l1_p1_col11_b = comp_l0_p2_col11_sum;
	
	assign u_comp_l1_p1_col11_cin = comp_l0_p2_col10_cout;
	
	assign u_comp_l1_p1_col12_a = comp_l0_p1_col11_cout;
	
	assign u_comp_l1_p1_col12_b = comp_l0_p2_col12_sum;
	
	assign u_comp_l1_p1_col12_cin = comp_l0_p2_col11_cout;
	
	assign u_comp_l1_p1_col13_a = comp_l0_p1_col12_cout;
	
	assign u_comp_l1_p1_col13_b = comp_l0_p2_col13_sum;
	
	assign u_comp_l1_p1_col13_cin = comp_l0_p2_col12_cout;
	
	assign u_comp_l1_p1_col14_a = comp_l0_p1_col13_cout;
	
	assign u_comp_l1_p1_col14_b = comp_l0_p2_col14_sum;
	
	assign u_comp_l1_p1_col14_cin = comp_l0_p2_col13_cout;
	
	assign u_comp_l1_p1_col15_a = comp_l0_p1_col14_cout;
	
	assign u_comp_l1_p1_col15_b = comp_l0_p2_col15_sum;
	
	assign u_comp_l1_p1_col15_cin = comp_l0_p2_col14_cout;
	
	assign u_comp_l1_p1_col16_a = comp_l0_p1_col15_cout;
	
	assign u_comp_l1_p1_col16_b = comp_l0_p2_col16_sum;
	
	assign u_comp_l1_p1_col16_cin = comp_l0_p2_col15_cout;
	
	assign u_comp_l1_p1_col17_a = comp_l0_p1_col16_cout;
	
	assign u_comp_l1_p1_col17_b = comp_l0_p2_col17_sum;
	
	assign u_comp_l1_p1_col17_cin = comp_l0_p2_col16_cout;
	
	assign u_comp_l1_p1_col18_a = comp_l0_p1_col17_cout;
	
	assign u_comp_l1_p1_col18_b = comp_l0_p2_col18_sum;
	
	assign u_comp_l1_p1_col18_cin = comp_l0_p2_col17_cout;
	
	assign u_comp_l1_p1_col19_a = comp_l0_p1_col18_cout;
	
	assign u_comp_l1_p1_col19_b = comp_l0_p2_col19_sum;
	
	assign u_comp_l1_p1_col19_cin = comp_l0_p2_col18_cout;
	
	assign u_comp_l1_p1_col20_a = comp_l0_p1_col19_cout;
	
	assign u_comp_l1_p1_col20_b = comp_l0_p2_col20_sum;
	
	assign u_comp_l1_p1_col20_cin = comp_l0_p2_col19_cout;
	
	assign u_comp_l1_p1_col21_a = comp_l0_p1_col20_cout;
	
	assign u_comp_l1_p1_col21_b = comp_l0_p2_col21_sum;
	
	assign u_comp_l1_p1_col21_cin = comp_l0_p2_col20_cout;
	
	assign u_comp_l1_p1_col22_a = comp_l0_p1_col21_cout;
	
	assign u_comp_l1_p1_col22_b = comp_l0_p2_col22_sum;
	
	assign u_comp_l1_p1_col22_cin = comp_l0_p2_col21_cout;
	
	assign u_comp_l1_p1_col23_a = comp_l0_p1_col22_cout;
	
	assign u_comp_l1_p1_col23_b = comp_l0_p2_col23_sum;
	
	assign u_comp_l1_p1_col23_cin = comp_l0_p2_col22_cout;
	
	assign u_comp_l1_p1_col24_a = comp_l0_p1_col23_cout;
	
	assign u_comp_l1_p1_col24_b = comp_l0_p2_col24_sum;
	
	assign u_comp_l1_p1_col24_cin = comp_l0_p2_col23_cout;
	
	assign u_comp_l1_p1_col25_a = comp_l0_p1_col24_cout;
	
	assign u_comp_l1_p1_col25_b = comp_l0_p2_col25_sum;
	
	assign u_comp_l1_p1_col25_cin = comp_l0_p2_col24_cout;
	
	assign u_comp_l1_p1_col26_a = comp_l0_p1_col25_cout;
	
	assign u_comp_l1_p1_col26_b = comp_l0_p2_col26_sum;
	
	assign u_comp_l1_p1_col26_cin = comp_l0_p2_col25_cout;
	
	assign u_comp_l1_p1_col27_a = comp_l0_p1_col26_cout;
	
	assign u_comp_l1_p1_col27_b = comp_l0_p2_col27_sum;
	
	assign u_comp_l1_p1_col27_cin = comp_l0_p2_col26_cout;
	
	assign u_comp_l1_p1_col28_a = comp_l0_p1_col27_cout;
	
	assign u_comp_l1_p1_col28_b = comp_l0_p2_col28_sum;
	
	assign u_comp_l1_p1_col28_cin = comp_l0_p2_col27_cout;
	
	assign u_comp_l1_p1_col29_a = comp_l0_p1_col28_cout;
	
	assign u_comp_l1_p1_col29_b = comp_l0_p2_col29_sum;
	
	assign u_comp_l1_p1_col29_cin = comp_l0_p2_col28_cout;
	
	assign u_comp_l1_p1_col30_a = comp_l0_p1_col29_cout;
	
	assign u_comp_l1_p1_col30_b = comp_l0_p2_col30_sum;
	
	assign u_comp_l1_p1_col30_cin = comp_l0_p2_col29_cout;
	
	assign u_comp_l1_p1_col31_a = comp_l0_p1_col30_cout;
	
	assign u_comp_l1_p1_col31_b = comp_l0_p2_col31_sum;
	
	assign u_comp_l1_p1_col31_cin = comp_l0_p2_col30_cout;
	
	assign u_comp_l2_p0_col0_a = comp_l1_p0_col0_sum;
	
	assign u_comp_l2_p0_col0_b = comp_pad_l1_p0;
	
	assign u_comp_l2_p0_col0_cin = comp_l1_p1_col0_sum;
	
	assign u_comp_l2_p0_col1_a = comp_l1_p0_col1_sum;
	
	assign u_comp_l2_p0_col1_b = comp_l1_p0_col0_cout;
	
	assign u_comp_l2_p0_col1_cin = comp_l1_p1_col1_sum;
	
	assign u_comp_l2_p0_col2_a = comp_l1_p0_col2_sum;
	
	assign u_comp_l2_p0_col2_b = comp_l1_p0_col1_cout;
	
	assign u_comp_l2_p0_col2_cin = comp_l1_p1_col2_sum;
	
	assign u_comp_l2_p0_col3_a = comp_l1_p0_col3_sum;
	
	assign u_comp_l2_p0_col3_b = comp_l1_p0_col2_cout;
	
	assign u_comp_l2_p0_col3_cin = comp_l1_p1_col3_sum;
	
	assign u_comp_l2_p0_col4_a = comp_l1_p0_col4_sum;
	
	assign u_comp_l2_p0_col4_b = comp_l1_p0_col3_cout;
	
	assign u_comp_l2_p0_col4_cin = comp_l1_p1_col4_sum;
	
	assign u_comp_l2_p0_col5_a = comp_l1_p0_col5_sum;
	
	assign u_comp_l2_p0_col5_b = comp_l1_p0_col4_cout;
	
	assign u_comp_l2_p0_col5_cin = comp_l1_p1_col5_sum;
	
	assign u_comp_l2_p0_col6_a = comp_l1_p0_col6_sum;
	
	assign u_comp_l2_p0_col6_b = comp_l1_p0_col5_cout;
	
	assign u_comp_l2_p0_col6_cin = comp_l1_p1_col6_sum;
	
	assign u_comp_l2_p0_col7_a = comp_l1_p0_col7_sum;
	
	assign u_comp_l2_p0_col7_b = comp_l1_p0_col6_cout;
	
	assign u_comp_l2_p0_col7_cin = comp_l1_p1_col7_sum;
	
	assign u_comp_l2_p0_col8_a = comp_l1_p0_col8_sum;
	
	assign u_comp_l2_p0_col8_b = comp_l1_p0_col7_cout;
	
	assign u_comp_l2_p0_col8_cin = comp_l1_p1_col8_sum;
	
	assign u_comp_l2_p0_col9_a = comp_l1_p0_col9_sum;
	
	assign u_comp_l2_p0_col9_b = comp_l1_p0_col8_cout;
	
	assign u_comp_l2_p0_col9_cin = comp_l1_p1_col9_sum;
	
	assign u_comp_l2_p0_col10_a = comp_l1_p0_col10_sum;
	
	assign u_comp_l2_p0_col10_b = comp_l1_p0_col9_cout;
	
	assign u_comp_l2_p0_col10_cin = comp_l1_p1_col10_sum;
	
	assign u_comp_l2_p0_col11_a = comp_l1_p0_col11_sum;
	
	assign u_comp_l2_p0_col11_b = comp_l1_p0_col10_cout;
	
	assign u_comp_l2_p0_col11_cin = comp_l1_p1_col11_sum;
	
	assign u_comp_l2_p0_col12_a = comp_l1_p0_col12_sum;
	
	assign u_comp_l2_p0_col12_b = comp_l1_p0_col11_cout;
	
	assign u_comp_l2_p0_col12_cin = comp_l1_p1_col12_sum;
	
	assign u_comp_l2_p0_col13_a = comp_l1_p0_col13_sum;
	
	assign u_comp_l2_p0_col13_b = comp_l1_p0_col12_cout;
	
	assign u_comp_l2_p0_col13_cin = comp_l1_p1_col13_sum;
	
	assign u_comp_l2_p0_col14_a = comp_l1_p0_col14_sum;
	
	assign u_comp_l2_p0_col14_b = comp_l1_p0_col13_cout;
	
	assign u_comp_l2_p0_col14_cin = comp_l1_p1_col14_sum;
	
	assign u_comp_l2_p0_col15_a = comp_l1_p0_col15_sum;
	
	assign u_comp_l2_p0_col15_b = comp_l1_p0_col14_cout;
	
	assign u_comp_l2_p0_col15_cin = comp_l1_p1_col15_sum;
	
	assign u_comp_l2_p0_col16_a = comp_l1_p0_col16_sum;
	
	assign u_comp_l2_p0_col16_b = comp_l1_p0_col15_cout;
	
	assign u_comp_l2_p0_col16_cin = comp_l1_p1_col16_sum;
	
	assign u_comp_l2_p0_col17_a = comp_l1_p0_col17_sum;
	
	assign u_comp_l2_p0_col17_b = comp_l1_p0_col16_cout;
	
	assign u_comp_l2_p0_col17_cin = comp_l1_p1_col17_sum;
	
	assign u_comp_l2_p0_col18_a = comp_l1_p0_col18_sum;
	
	assign u_comp_l2_p0_col18_b = comp_l1_p0_col17_cout;
	
	assign u_comp_l2_p0_col18_cin = comp_l1_p1_col18_sum;
	
	assign u_comp_l2_p0_col19_a = comp_l1_p0_col19_sum;
	
	assign u_comp_l2_p0_col19_b = comp_l1_p0_col18_cout;
	
	assign u_comp_l2_p0_col19_cin = comp_l1_p1_col19_sum;
	
	assign u_comp_l2_p0_col20_a = comp_l1_p0_col20_sum;
	
	assign u_comp_l2_p0_col20_b = comp_l1_p0_col19_cout;
	
	assign u_comp_l2_p0_col20_cin = comp_l1_p1_col20_sum;
	
	assign u_comp_l2_p0_col21_a = comp_l1_p0_col21_sum;
	
	assign u_comp_l2_p0_col21_b = comp_l1_p0_col20_cout;
	
	assign u_comp_l2_p0_col21_cin = comp_l1_p1_col21_sum;
	
	assign u_comp_l2_p0_col22_a = comp_l1_p0_col22_sum;
	
	assign u_comp_l2_p0_col22_b = comp_l1_p0_col21_cout;
	
	assign u_comp_l2_p0_col22_cin = comp_l1_p1_col22_sum;
	
	assign u_comp_l2_p0_col23_a = comp_l1_p0_col23_sum;
	
	assign u_comp_l2_p0_col23_b = comp_l1_p0_col22_cout;
	
	assign u_comp_l2_p0_col23_cin = comp_l1_p1_col23_sum;
	
	assign u_comp_l2_p0_col24_a = comp_l1_p0_col24_sum;
	
	assign u_comp_l2_p0_col24_b = comp_l1_p0_col23_cout;
	
	assign u_comp_l2_p0_col24_cin = comp_l1_p1_col24_sum;
	
	assign u_comp_l2_p0_col25_a = comp_l1_p0_col25_sum;
	
	assign u_comp_l2_p0_col25_b = comp_l1_p0_col24_cout;
	
	assign u_comp_l2_p0_col25_cin = comp_l1_p1_col25_sum;
	
	assign u_comp_l2_p0_col26_a = comp_l1_p0_col26_sum;
	
	assign u_comp_l2_p0_col26_b = comp_l1_p0_col25_cout;
	
	assign u_comp_l2_p0_col26_cin = comp_l1_p1_col26_sum;
	
	assign u_comp_l2_p0_col27_a = comp_l1_p0_col27_sum;
	
	assign u_comp_l2_p0_col27_b = comp_l1_p0_col26_cout;
	
	assign u_comp_l2_p0_col27_cin = comp_l1_p1_col27_sum;
	
	assign u_comp_l2_p0_col28_a = comp_l1_p0_col28_sum;
	
	assign u_comp_l2_p0_col28_b = comp_l1_p0_col27_cout;
	
	assign u_comp_l2_p0_col28_cin = comp_l1_p1_col28_sum;
	
	assign u_comp_l2_p0_col29_a = comp_l1_p0_col29_sum;
	
	assign u_comp_l2_p0_col29_b = comp_l1_p0_col28_cout;
	
	assign u_comp_l2_p0_col29_cin = comp_l1_p1_col29_sum;
	
	assign u_comp_l2_p0_col30_a = comp_l1_p0_col30_sum;
	
	assign u_comp_l2_p0_col30_b = comp_l1_p0_col29_cout;
	
	assign u_comp_l2_p0_col30_cin = comp_l1_p1_col30_sum;
	
	assign u_comp_l2_p0_col31_a = comp_l1_p0_col31_sum;
	
	assign u_comp_l2_p0_col31_b = comp_l1_p0_col30_cout;
	
	assign u_comp_l2_p0_col31_cin = comp_l1_p1_col31_sum;
	
	assign u_comp_l3_p0_col0_a = comp_l2_p0_col0_sum;
	
	assign u_comp_l3_p0_col0_b = comp_pad_l2_p0;
	
	assign u_comp_l3_p0_col0_cin = comp_pad_l1_p1;
	
	assign u_comp_l3_p0_col1_a = comp_l2_p0_col1_sum;
	
	assign u_comp_l3_p0_col1_b = comp_l2_p0_col0_cout;
	
	assign u_comp_l3_p0_col1_cin = comp_l1_p1_col0_cout;
	
	assign u_comp_l3_p0_col2_a = comp_l2_p0_col2_sum;
	
	assign u_comp_l3_p0_col2_b = comp_l2_p0_col1_cout;
	
	assign u_comp_l3_p0_col2_cin = comp_l1_p1_col1_cout;
	
	assign u_comp_l3_p0_col3_a = comp_l2_p0_col3_sum;
	
	assign u_comp_l3_p0_col3_b = comp_l2_p0_col2_cout;
	
	assign u_comp_l3_p0_col3_cin = comp_l1_p1_col2_cout;
	
	assign u_comp_l3_p0_col4_a = comp_l2_p0_col4_sum;
	
	assign u_comp_l3_p0_col4_b = comp_l2_p0_col3_cout;
	
	assign u_comp_l3_p0_col4_cin = comp_l1_p1_col3_cout;
	
	assign u_comp_l3_p0_col5_a = comp_l2_p0_col5_sum;
	
	assign u_comp_l3_p0_col5_b = comp_l2_p0_col4_cout;
	
	assign u_comp_l3_p0_col5_cin = comp_l1_p1_col4_cout;
	
	assign u_comp_l3_p0_col6_a = comp_l2_p0_col6_sum;
	
	assign u_comp_l3_p0_col6_b = comp_l2_p0_col5_cout;
	
	assign u_comp_l3_p0_col6_cin = comp_l1_p1_col5_cout;
	
	assign u_comp_l3_p0_col7_a = comp_l2_p0_col7_sum;
	
	assign u_comp_l3_p0_col7_b = comp_l2_p0_col6_cout;
	
	assign u_comp_l3_p0_col7_cin = comp_l1_p1_col6_cout;
	
	assign u_comp_l3_p0_col8_a = comp_l2_p0_col8_sum;
	
	assign u_comp_l3_p0_col8_b = comp_l2_p0_col7_cout;
	
	assign u_comp_l3_p0_col8_cin = comp_l1_p1_col7_cout;
	
	assign u_comp_l3_p0_col9_a = comp_l2_p0_col9_sum;
	
	assign u_comp_l3_p0_col9_b = comp_l2_p0_col8_cout;
	
	assign u_comp_l3_p0_col9_cin = comp_l1_p1_col8_cout;
	
	assign u_comp_l3_p0_col10_a = comp_l2_p0_col10_sum;
	
	assign u_comp_l3_p0_col10_b = comp_l2_p0_col9_cout;
	
	assign u_comp_l3_p0_col10_cin = comp_l1_p1_col9_cout;
	
	assign u_comp_l3_p0_col11_a = comp_l2_p0_col11_sum;
	
	assign u_comp_l3_p0_col11_b = comp_l2_p0_col10_cout;
	
	assign u_comp_l3_p0_col11_cin = comp_l1_p1_col10_cout;
	
	assign u_comp_l3_p0_col12_a = comp_l2_p0_col12_sum;
	
	assign u_comp_l3_p0_col12_b = comp_l2_p0_col11_cout;
	
	assign u_comp_l3_p0_col12_cin = comp_l1_p1_col11_cout;
	
	assign u_comp_l3_p0_col13_a = comp_l2_p0_col13_sum;
	
	assign u_comp_l3_p0_col13_b = comp_l2_p0_col12_cout;
	
	assign u_comp_l3_p0_col13_cin = comp_l1_p1_col12_cout;
	
	assign u_comp_l3_p0_col14_a = comp_l2_p0_col14_sum;
	
	assign u_comp_l3_p0_col14_b = comp_l2_p0_col13_cout;
	
	assign u_comp_l3_p0_col14_cin = comp_l1_p1_col13_cout;
	
	assign u_comp_l3_p0_col15_a = comp_l2_p0_col15_sum;
	
	assign u_comp_l3_p0_col15_b = comp_l2_p0_col14_cout;
	
	assign u_comp_l3_p0_col15_cin = comp_l1_p1_col14_cout;
	
	assign u_comp_l3_p0_col16_a = comp_l2_p0_col16_sum;
	
	assign u_comp_l3_p0_col16_b = comp_l2_p0_col15_cout;
	
	assign u_comp_l3_p0_col16_cin = comp_l1_p1_col15_cout;
	
	assign u_comp_l3_p0_col17_a = comp_l2_p0_col17_sum;
	
	assign u_comp_l3_p0_col17_b = comp_l2_p0_col16_cout;
	
	assign u_comp_l3_p0_col17_cin = comp_l1_p1_col16_cout;
	
	assign u_comp_l3_p0_col18_a = comp_l2_p0_col18_sum;
	
	assign u_comp_l3_p0_col18_b = comp_l2_p0_col17_cout;
	
	assign u_comp_l3_p0_col18_cin = comp_l1_p1_col17_cout;
	
	assign u_comp_l3_p0_col19_a = comp_l2_p0_col19_sum;
	
	assign u_comp_l3_p0_col19_b = comp_l2_p0_col18_cout;
	
	assign u_comp_l3_p0_col19_cin = comp_l1_p1_col18_cout;
	
	assign u_comp_l3_p0_col20_a = comp_l2_p0_col20_sum;
	
	assign u_comp_l3_p0_col20_b = comp_l2_p0_col19_cout;
	
	assign u_comp_l3_p0_col20_cin = comp_l1_p1_col19_cout;
	
	assign u_comp_l3_p0_col21_a = comp_l2_p0_col21_sum;
	
	assign u_comp_l3_p0_col21_b = comp_l2_p0_col20_cout;
	
	assign u_comp_l3_p0_col21_cin = comp_l1_p1_col20_cout;
	
	assign u_comp_l3_p0_col22_a = comp_l2_p0_col22_sum;
	
	assign u_comp_l3_p0_col22_b = comp_l2_p0_col21_cout;
	
	assign u_comp_l3_p0_col22_cin = comp_l1_p1_col21_cout;
	
	assign u_comp_l3_p0_col23_a = comp_l2_p0_col23_sum;
	
	assign u_comp_l3_p0_col23_b = comp_l2_p0_col22_cout;
	
	assign u_comp_l3_p0_col23_cin = comp_l1_p1_col22_cout;
	
	assign u_comp_l3_p0_col24_a = comp_l2_p0_col24_sum;
	
	assign u_comp_l3_p0_col24_b = comp_l2_p0_col23_cout;
	
	assign u_comp_l3_p0_col24_cin = comp_l1_p1_col23_cout;
	
	assign u_comp_l3_p0_col25_a = comp_l2_p0_col25_sum;
	
	assign u_comp_l3_p0_col25_b = comp_l2_p0_col24_cout;
	
	assign u_comp_l3_p0_col25_cin = comp_l1_p1_col24_cout;
	
	assign u_comp_l3_p0_col26_a = comp_l2_p0_col26_sum;
	
	assign u_comp_l3_p0_col26_b = comp_l2_p0_col25_cout;
	
	assign u_comp_l3_p0_col26_cin = comp_l1_p1_col25_cout;
	
	assign u_comp_l3_p0_col27_a = comp_l2_p0_col27_sum;
	
	assign u_comp_l3_p0_col27_b = comp_l2_p0_col26_cout;
	
	assign u_comp_l3_p0_col27_cin = comp_l1_p1_col26_cout;
	
	assign u_comp_l3_p0_col28_a = comp_l2_p0_col28_sum;
	
	assign u_comp_l3_p0_col28_b = comp_l2_p0_col27_cout;
	
	assign u_comp_l3_p0_col28_cin = comp_l1_p1_col27_cout;
	
	assign u_comp_l3_p0_col29_a = comp_l2_p0_col29_sum;
	
	assign u_comp_l3_p0_col29_b = comp_l2_p0_col28_cout;
	
	assign u_comp_l3_p0_col29_cin = comp_l1_p1_col28_cout;
	
	assign u_comp_l3_p0_col30_a = comp_l2_p0_col30_sum;
	
	assign u_comp_l3_p0_col30_b = comp_l2_p0_col29_cout;
	
	assign u_comp_l3_p0_col30_cin = comp_l1_p1_col29_cout;
	
	assign u_comp_l3_p0_col31_a = comp_l2_p0_col31_sum;
	
	assign u_comp_l3_p0_col31_b = comp_l2_p0_col30_cout;
	
	assign u_comp_l3_p0_col31_cin = comp_l1_p1_col30_cout;
	
	assign u_comp_l4_p0_col0_a = comp_l3_p0_col0_sum;
	
	assign u_comp_l4_p0_col0_b = comp_pad_l3_p0;
	
	assign u_comp_l4_p0_col0_cin = p_9_0;
	
	assign u_comp_l4_p0_col1_a = comp_l3_p0_col1_sum;
	
	assign u_comp_l4_p0_col1_b = comp_l3_p0_col0_cout;
	
	assign u_comp_l4_p0_col1_cin = p_9_1;
	
	assign u_comp_l4_p0_col2_a = comp_l3_p0_col2_sum;
	
	assign u_comp_l4_p0_col2_b = comp_l3_p0_col1_cout;
	
	assign u_comp_l4_p0_col2_cin = p_9_2;
	
	assign u_comp_l4_p0_col3_a = comp_l3_p0_col3_sum;
	
	assign u_comp_l4_p0_col3_b = comp_l3_p0_col2_cout;
	
	assign u_comp_l4_p0_col3_cin = p_9_3;
	
	assign u_comp_l4_p0_col4_a = comp_l3_p0_col4_sum;
	
	assign u_comp_l4_p0_col4_b = comp_l3_p0_col3_cout;
	
	assign u_comp_l4_p0_col4_cin = p_9_4;
	
	assign u_comp_l4_p0_col5_a = comp_l3_p0_col5_sum;
	
	assign u_comp_l4_p0_col5_b = comp_l3_p0_col4_cout;
	
	assign u_comp_l4_p0_col5_cin = p_9_5;
	
	assign u_comp_l4_p0_col6_a = comp_l3_p0_col6_sum;
	
	assign u_comp_l4_p0_col6_b = comp_l3_p0_col5_cout;
	
	assign u_comp_l4_p0_col6_cin = p_9_6;
	
	assign u_comp_l4_p0_col7_a = comp_l3_p0_col7_sum;
	
	assign u_comp_l4_p0_col7_b = comp_l3_p0_col6_cout;
	
	assign u_comp_l4_p0_col7_cin = p_9_7;
	
	assign u_comp_l4_p0_col8_a = comp_l3_p0_col8_sum;
	
	assign u_comp_l4_p0_col8_b = comp_l3_p0_col7_cout;
	
	assign u_comp_l4_p0_col8_cin = p_9_8;
	
	assign u_comp_l4_p0_col9_a = comp_l3_p0_col9_sum;
	
	assign u_comp_l4_p0_col9_b = comp_l3_p0_col8_cout;
	
	assign u_comp_l4_p0_col9_cin = p_9_9;
	
	assign u_comp_l4_p0_col10_a = comp_l3_p0_col10_sum;
	
	assign u_comp_l4_p0_col10_b = comp_l3_p0_col9_cout;
	
	assign u_comp_l4_p0_col10_cin = p_9_10;
	
	assign u_comp_l4_p0_col11_a = comp_l3_p0_col11_sum;
	
	assign u_comp_l4_p0_col11_b = comp_l3_p0_col10_cout;
	
	assign u_comp_l4_p0_col11_cin = p_9_11;
	
	assign u_comp_l4_p0_col12_a = comp_l3_p0_col12_sum;
	
	assign u_comp_l4_p0_col12_b = comp_l3_p0_col11_cout;
	
	assign u_comp_l4_p0_col12_cin = p_9_12;
	
	assign u_comp_l4_p0_col13_a = comp_l3_p0_col13_sum;
	
	assign u_comp_l4_p0_col13_b = comp_l3_p0_col12_cout;
	
	assign u_comp_l4_p0_col13_cin = p_9_13;
	
	assign u_comp_l4_p0_col14_a = comp_l3_p0_col14_sum;
	
	assign u_comp_l4_p0_col14_b = comp_l3_p0_col13_cout;
	
	assign u_comp_l4_p0_col14_cin = p_9_14;
	
	assign u_comp_l4_p0_col15_a = comp_l3_p0_col15_sum;
	
	assign u_comp_l4_p0_col15_b = comp_l3_p0_col14_cout;
	
	assign u_comp_l4_p0_col15_cin = p_9_15;
	
	assign u_comp_l4_p0_col16_a = comp_l3_p0_col16_sum;
	
	assign u_comp_l4_p0_col16_b = comp_l3_p0_col15_cout;
	
	assign u_comp_l4_p0_col16_cin = p_9_16;
	
	assign u_comp_l4_p0_col17_a = comp_l3_p0_col17_sum;
	
	assign u_comp_l4_p0_col17_b = comp_l3_p0_col16_cout;
	
	assign u_comp_l4_p0_col17_cin = p_9_17;
	
	assign u_comp_l4_p0_col18_a = comp_l3_p0_col18_sum;
	
	assign u_comp_l4_p0_col18_b = comp_l3_p0_col17_cout;
	
	assign u_comp_l4_p0_col18_cin = p_9_18;
	
	assign u_comp_l4_p0_col19_a = comp_l3_p0_col19_sum;
	
	assign u_comp_l4_p0_col19_b = comp_l3_p0_col18_cout;
	
	assign u_comp_l4_p0_col19_cin = p_9_19;
	
	assign u_comp_l4_p0_col20_a = comp_l3_p0_col20_sum;
	
	assign u_comp_l4_p0_col20_b = comp_l3_p0_col19_cout;
	
	assign u_comp_l4_p0_col20_cin = p_9_20;
	
	assign u_comp_l4_p0_col21_a = comp_l3_p0_col21_sum;
	
	assign u_comp_l4_p0_col21_b = comp_l3_p0_col20_cout;
	
	assign u_comp_l4_p0_col21_cin = p_9_21;
	
	assign u_comp_l4_p0_col22_a = comp_l3_p0_col22_sum;
	
	assign u_comp_l4_p0_col22_b = comp_l3_p0_col21_cout;
	
	assign u_comp_l4_p0_col22_cin = p_9_22;
	
	assign u_comp_l4_p0_col23_a = comp_l3_p0_col23_sum;
	
	assign u_comp_l4_p0_col23_b = comp_l3_p0_col22_cout;
	
	assign u_comp_l4_p0_col23_cin = p_9_23;
	
	assign u_comp_l4_p0_col24_a = comp_l3_p0_col24_sum;
	
	assign u_comp_l4_p0_col24_b = comp_l3_p0_col23_cout;
	
	assign u_comp_l4_p0_col24_cin = p_9_24;
	
	assign u_comp_l4_p0_col25_a = comp_l3_p0_col25_sum;
	
	assign u_comp_l4_p0_col25_b = comp_l3_p0_col24_cout;
	
	assign u_comp_l4_p0_col25_cin = p_9_25;
	
	assign u_comp_l4_p0_col26_a = comp_l3_p0_col26_sum;
	
	assign u_comp_l4_p0_col26_b = comp_l3_p0_col25_cout;
	
	assign u_comp_l4_p0_col26_cin = p_9_26;
	
	assign u_comp_l4_p0_col27_a = comp_l3_p0_col27_sum;
	
	assign u_comp_l4_p0_col27_b = comp_l3_p0_col26_cout;
	
	assign u_comp_l4_p0_col27_cin = p_9_27;
	
	assign u_comp_l4_p0_col28_a = comp_l3_p0_col28_sum;
	
	assign u_comp_l4_p0_col28_b = comp_l3_p0_col27_cout;
	
	assign u_comp_l4_p0_col28_cin = p_9_28;
	
	assign u_comp_l4_p0_col29_a = comp_l3_p0_col29_sum;
	
	assign u_comp_l4_p0_col29_b = comp_l3_p0_col28_cout;
	
	assign u_comp_l4_p0_col29_cin = p_9_29;
	
	assign u_comp_l4_p0_col30_a = comp_l3_p0_col30_sum;
	
	assign u_comp_l4_p0_col30_b = comp_l3_p0_col29_cout;
	
	assign u_comp_l4_p0_col30_cin = p_9_30;
	
	assign u_comp_l4_p0_col31_a = comp_l3_p0_col31_sum;
	
	assign u_comp_l4_p0_col31_b = comp_l3_p0_col30_cout;
	
	assign u_comp_l4_p0_col31_cin = p_9_31;
	

	//module inst.
	FullAdder u_comp_l0_p0_col0 (
		.a(u_comp_l0_p0_col0_a),
		.b(u_comp_l0_p0_col0_b),
		.cin(u_comp_l0_p0_col0_cin),
		.cout(u_comp_l0_p0_col0_cout),
		.sum(u_comp_l0_p0_col0_sum));
	FullAdder u_comp_l0_p0_col1 (
		.a(u_comp_l0_p0_col1_a),
		.b(u_comp_l0_p0_col1_b),
		.cin(u_comp_l0_p0_col1_cin),
		.cout(u_comp_l0_p0_col1_cout),
		.sum(u_comp_l0_p0_col1_sum));
	FullAdder u_comp_l0_p0_col2 (
		.a(u_comp_l0_p0_col2_a),
		.b(u_comp_l0_p0_col2_b),
		.cin(u_comp_l0_p0_col2_cin),
		.cout(u_comp_l0_p0_col2_cout),
		.sum(u_comp_l0_p0_col2_sum));
	FullAdder u_comp_l0_p0_col3 (
		.a(u_comp_l0_p0_col3_a),
		.b(u_comp_l0_p0_col3_b),
		.cin(u_comp_l0_p0_col3_cin),
		.cout(u_comp_l0_p0_col3_cout),
		.sum(u_comp_l0_p0_col3_sum));
	FullAdder u_comp_l0_p0_col4 (
		.a(u_comp_l0_p0_col4_a),
		.b(u_comp_l0_p0_col4_b),
		.cin(u_comp_l0_p0_col4_cin),
		.cout(u_comp_l0_p0_col4_cout),
		.sum(u_comp_l0_p0_col4_sum));
	FullAdder u_comp_l0_p0_col5 (
		.a(u_comp_l0_p0_col5_a),
		.b(u_comp_l0_p0_col5_b),
		.cin(u_comp_l0_p0_col5_cin),
		.cout(u_comp_l0_p0_col5_cout),
		.sum(u_comp_l0_p0_col5_sum));
	FullAdder u_comp_l0_p0_col6 (
		.a(u_comp_l0_p0_col6_a),
		.b(u_comp_l0_p0_col6_b),
		.cin(u_comp_l0_p0_col6_cin),
		.cout(u_comp_l0_p0_col6_cout),
		.sum(u_comp_l0_p0_col6_sum));
	FullAdder u_comp_l0_p0_col7 (
		.a(u_comp_l0_p0_col7_a),
		.b(u_comp_l0_p0_col7_b),
		.cin(u_comp_l0_p0_col7_cin),
		.cout(u_comp_l0_p0_col7_cout),
		.sum(u_comp_l0_p0_col7_sum));
	FullAdder u_comp_l0_p0_col8 (
		.a(u_comp_l0_p0_col8_a),
		.b(u_comp_l0_p0_col8_b),
		.cin(u_comp_l0_p0_col8_cin),
		.cout(u_comp_l0_p0_col8_cout),
		.sum(u_comp_l0_p0_col8_sum));
	FullAdder u_comp_l0_p0_col9 (
		.a(u_comp_l0_p0_col9_a),
		.b(u_comp_l0_p0_col9_b),
		.cin(u_comp_l0_p0_col9_cin),
		.cout(u_comp_l0_p0_col9_cout),
		.sum(u_comp_l0_p0_col9_sum));
	FullAdder u_comp_l0_p0_col10 (
		.a(u_comp_l0_p0_col10_a),
		.b(u_comp_l0_p0_col10_b),
		.cin(u_comp_l0_p0_col10_cin),
		.cout(u_comp_l0_p0_col10_cout),
		.sum(u_comp_l0_p0_col10_sum));
	FullAdder u_comp_l0_p0_col11 (
		.a(u_comp_l0_p0_col11_a),
		.b(u_comp_l0_p0_col11_b),
		.cin(u_comp_l0_p0_col11_cin),
		.cout(u_comp_l0_p0_col11_cout),
		.sum(u_comp_l0_p0_col11_sum));
	FullAdder u_comp_l0_p0_col12 (
		.a(u_comp_l0_p0_col12_a),
		.b(u_comp_l0_p0_col12_b),
		.cin(u_comp_l0_p0_col12_cin),
		.cout(u_comp_l0_p0_col12_cout),
		.sum(u_comp_l0_p0_col12_sum));
	FullAdder u_comp_l0_p0_col13 (
		.a(u_comp_l0_p0_col13_a),
		.b(u_comp_l0_p0_col13_b),
		.cin(u_comp_l0_p0_col13_cin),
		.cout(u_comp_l0_p0_col13_cout),
		.sum(u_comp_l0_p0_col13_sum));
	FullAdder u_comp_l0_p0_col14 (
		.a(u_comp_l0_p0_col14_a),
		.b(u_comp_l0_p0_col14_b),
		.cin(u_comp_l0_p0_col14_cin),
		.cout(u_comp_l0_p0_col14_cout),
		.sum(u_comp_l0_p0_col14_sum));
	FullAdder u_comp_l0_p0_col15 (
		.a(u_comp_l0_p0_col15_a),
		.b(u_comp_l0_p0_col15_b),
		.cin(u_comp_l0_p0_col15_cin),
		.cout(u_comp_l0_p0_col15_cout),
		.sum(u_comp_l0_p0_col15_sum));
	FullAdder u_comp_l0_p0_col16 (
		.a(u_comp_l0_p0_col16_a),
		.b(u_comp_l0_p0_col16_b),
		.cin(u_comp_l0_p0_col16_cin),
		.cout(u_comp_l0_p0_col16_cout),
		.sum(u_comp_l0_p0_col16_sum));
	FullAdder u_comp_l0_p0_col17 (
		.a(u_comp_l0_p0_col17_a),
		.b(u_comp_l0_p0_col17_b),
		.cin(u_comp_l0_p0_col17_cin),
		.cout(u_comp_l0_p0_col17_cout),
		.sum(u_comp_l0_p0_col17_sum));
	FullAdder u_comp_l0_p0_col18 (
		.a(u_comp_l0_p0_col18_a),
		.b(u_comp_l0_p0_col18_b),
		.cin(u_comp_l0_p0_col18_cin),
		.cout(u_comp_l0_p0_col18_cout),
		.sum(u_comp_l0_p0_col18_sum));
	FullAdder u_comp_l0_p0_col19 (
		.a(u_comp_l0_p0_col19_a),
		.b(u_comp_l0_p0_col19_b),
		.cin(u_comp_l0_p0_col19_cin),
		.cout(u_comp_l0_p0_col19_cout),
		.sum(u_comp_l0_p0_col19_sum));
	FullAdder u_comp_l0_p0_col20 (
		.a(u_comp_l0_p0_col20_a),
		.b(u_comp_l0_p0_col20_b),
		.cin(u_comp_l0_p0_col20_cin),
		.cout(u_comp_l0_p0_col20_cout),
		.sum(u_comp_l0_p0_col20_sum));
	FullAdder u_comp_l0_p0_col21 (
		.a(u_comp_l0_p0_col21_a),
		.b(u_comp_l0_p0_col21_b),
		.cin(u_comp_l0_p0_col21_cin),
		.cout(u_comp_l0_p0_col21_cout),
		.sum(u_comp_l0_p0_col21_sum));
	FullAdder u_comp_l0_p0_col22 (
		.a(u_comp_l0_p0_col22_a),
		.b(u_comp_l0_p0_col22_b),
		.cin(u_comp_l0_p0_col22_cin),
		.cout(u_comp_l0_p0_col22_cout),
		.sum(u_comp_l0_p0_col22_sum));
	FullAdder u_comp_l0_p0_col23 (
		.a(u_comp_l0_p0_col23_a),
		.b(u_comp_l0_p0_col23_b),
		.cin(u_comp_l0_p0_col23_cin),
		.cout(u_comp_l0_p0_col23_cout),
		.sum(u_comp_l0_p0_col23_sum));
	FullAdder u_comp_l0_p0_col24 (
		.a(u_comp_l0_p0_col24_a),
		.b(u_comp_l0_p0_col24_b),
		.cin(u_comp_l0_p0_col24_cin),
		.cout(u_comp_l0_p0_col24_cout),
		.sum(u_comp_l0_p0_col24_sum));
	FullAdder u_comp_l0_p0_col25 (
		.a(u_comp_l0_p0_col25_a),
		.b(u_comp_l0_p0_col25_b),
		.cin(u_comp_l0_p0_col25_cin),
		.cout(u_comp_l0_p0_col25_cout),
		.sum(u_comp_l0_p0_col25_sum));
	FullAdder u_comp_l0_p0_col26 (
		.a(u_comp_l0_p0_col26_a),
		.b(u_comp_l0_p0_col26_b),
		.cin(u_comp_l0_p0_col26_cin),
		.cout(u_comp_l0_p0_col26_cout),
		.sum(u_comp_l0_p0_col26_sum));
	FullAdder u_comp_l0_p0_col27 (
		.a(u_comp_l0_p0_col27_a),
		.b(u_comp_l0_p0_col27_b),
		.cin(u_comp_l0_p0_col27_cin),
		.cout(u_comp_l0_p0_col27_cout),
		.sum(u_comp_l0_p0_col27_sum));
	FullAdder u_comp_l0_p0_col28 (
		.a(u_comp_l0_p0_col28_a),
		.b(u_comp_l0_p0_col28_b),
		.cin(u_comp_l0_p0_col28_cin),
		.cout(u_comp_l0_p0_col28_cout),
		.sum(u_comp_l0_p0_col28_sum));
	FullAdder u_comp_l0_p0_col29 (
		.a(u_comp_l0_p0_col29_a),
		.b(u_comp_l0_p0_col29_b),
		.cin(u_comp_l0_p0_col29_cin),
		.cout(u_comp_l0_p0_col29_cout),
		.sum(u_comp_l0_p0_col29_sum));
	FullAdder u_comp_l0_p0_col30 (
		.a(u_comp_l0_p0_col30_a),
		.b(u_comp_l0_p0_col30_b),
		.cin(u_comp_l0_p0_col30_cin),
		.cout(u_comp_l0_p0_col30_cout),
		.sum(u_comp_l0_p0_col30_sum));
	FullAdder u_comp_l0_p0_col31 (
		.a(u_comp_l0_p0_col31_a),
		.b(u_comp_l0_p0_col31_b),
		.cin(u_comp_l0_p0_col31_cin),
		.cout(comp_l0_p0_col31_cout),
		.sum(u_comp_l0_p0_col31_sum));
	FullAdder u_comp_l0_p1_col0 (
		.a(u_comp_l0_p1_col0_a),
		.b(u_comp_l0_p1_col0_b),
		.cin(u_comp_l0_p1_col0_cin),
		.cout(u_comp_l0_p1_col0_cout),
		.sum(u_comp_l0_p1_col0_sum));
	FullAdder u_comp_l0_p1_col1 (
		.a(u_comp_l0_p1_col1_a),
		.b(u_comp_l0_p1_col1_b),
		.cin(u_comp_l0_p1_col1_cin),
		.cout(u_comp_l0_p1_col1_cout),
		.sum(u_comp_l0_p1_col1_sum));
	FullAdder u_comp_l0_p1_col2 (
		.a(u_comp_l0_p1_col2_a),
		.b(u_comp_l0_p1_col2_b),
		.cin(u_comp_l0_p1_col2_cin),
		.cout(u_comp_l0_p1_col2_cout),
		.sum(u_comp_l0_p1_col2_sum));
	FullAdder u_comp_l0_p1_col3 (
		.a(u_comp_l0_p1_col3_a),
		.b(u_comp_l0_p1_col3_b),
		.cin(u_comp_l0_p1_col3_cin),
		.cout(u_comp_l0_p1_col3_cout),
		.sum(u_comp_l0_p1_col3_sum));
	FullAdder u_comp_l0_p1_col4 (
		.a(u_comp_l0_p1_col4_a),
		.b(u_comp_l0_p1_col4_b),
		.cin(u_comp_l0_p1_col4_cin),
		.cout(u_comp_l0_p1_col4_cout),
		.sum(u_comp_l0_p1_col4_sum));
	FullAdder u_comp_l0_p1_col5 (
		.a(u_comp_l0_p1_col5_a),
		.b(u_comp_l0_p1_col5_b),
		.cin(u_comp_l0_p1_col5_cin),
		.cout(u_comp_l0_p1_col5_cout),
		.sum(u_comp_l0_p1_col5_sum));
	FullAdder u_comp_l0_p1_col6 (
		.a(u_comp_l0_p1_col6_a),
		.b(u_comp_l0_p1_col6_b),
		.cin(u_comp_l0_p1_col6_cin),
		.cout(u_comp_l0_p1_col6_cout),
		.sum(u_comp_l0_p1_col6_sum));
	FullAdder u_comp_l0_p1_col7 (
		.a(u_comp_l0_p1_col7_a),
		.b(u_comp_l0_p1_col7_b),
		.cin(u_comp_l0_p1_col7_cin),
		.cout(u_comp_l0_p1_col7_cout),
		.sum(u_comp_l0_p1_col7_sum));
	FullAdder u_comp_l0_p1_col8 (
		.a(u_comp_l0_p1_col8_a),
		.b(u_comp_l0_p1_col8_b),
		.cin(u_comp_l0_p1_col8_cin),
		.cout(u_comp_l0_p1_col8_cout),
		.sum(u_comp_l0_p1_col8_sum));
	FullAdder u_comp_l0_p1_col9 (
		.a(u_comp_l0_p1_col9_a),
		.b(u_comp_l0_p1_col9_b),
		.cin(u_comp_l0_p1_col9_cin),
		.cout(u_comp_l0_p1_col9_cout),
		.sum(u_comp_l0_p1_col9_sum));
	FullAdder u_comp_l0_p1_col10 (
		.a(u_comp_l0_p1_col10_a),
		.b(u_comp_l0_p1_col10_b),
		.cin(u_comp_l0_p1_col10_cin),
		.cout(u_comp_l0_p1_col10_cout),
		.sum(u_comp_l0_p1_col10_sum));
	FullAdder u_comp_l0_p1_col11 (
		.a(u_comp_l0_p1_col11_a),
		.b(u_comp_l0_p1_col11_b),
		.cin(u_comp_l0_p1_col11_cin),
		.cout(u_comp_l0_p1_col11_cout),
		.sum(u_comp_l0_p1_col11_sum));
	FullAdder u_comp_l0_p1_col12 (
		.a(u_comp_l0_p1_col12_a),
		.b(u_comp_l0_p1_col12_b),
		.cin(u_comp_l0_p1_col12_cin),
		.cout(u_comp_l0_p1_col12_cout),
		.sum(u_comp_l0_p1_col12_sum));
	FullAdder u_comp_l0_p1_col13 (
		.a(u_comp_l0_p1_col13_a),
		.b(u_comp_l0_p1_col13_b),
		.cin(u_comp_l0_p1_col13_cin),
		.cout(u_comp_l0_p1_col13_cout),
		.sum(u_comp_l0_p1_col13_sum));
	FullAdder u_comp_l0_p1_col14 (
		.a(u_comp_l0_p1_col14_a),
		.b(u_comp_l0_p1_col14_b),
		.cin(u_comp_l0_p1_col14_cin),
		.cout(u_comp_l0_p1_col14_cout),
		.sum(u_comp_l0_p1_col14_sum));
	FullAdder u_comp_l0_p1_col15 (
		.a(u_comp_l0_p1_col15_a),
		.b(u_comp_l0_p1_col15_b),
		.cin(u_comp_l0_p1_col15_cin),
		.cout(u_comp_l0_p1_col15_cout),
		.sum(u_comp_l0_p1_col15_sum));
	FullAdder u_comp_l0_p1_col16 (
		.a(u_comp_l0_p1_col16_a),
		.b(u_comp_l0_p1_col16_b),
		.cin(u_comp_l0_p1_col16_cin),
		.cout(u_comp_l0_p1_col16_cout),
		.sum(u_comp_l0_p1_col16_sum));
	FullAdder u_comp_l0_p1_col17 (
		.a(u_comp_l0_p1_col17_a),
		.b(u_comp_l0_p1_col17_b),
		.cin(u_comp_l0_p1_col17_cin),
		.cout(u_comp_l0_p1_col17_cout),
		.sum(u_comp_l0_p1_col17_sum));
	FullAdder u_comp_l0_p1_col18 (
		.a(u_comp_l0_p1_col18_a),
		.b(u_comp_l0_p1_col18_b),
		.cin(u_comp_l0_p1_col18_cin),
		.cout(u_comp_l0_p1_col18_cout),
		.sum(u_comp_l0_p1_col18_sum));
	FullAdder u_comp_l0_p1_col19 (
		.a(u_comp_l0_p1_col19_a),
		.b(u_comp_l0_p1_col19_b),
		.cin(u_comp_l0_p1_col19_cin),
		.cout(u_comp_l0_p1_col19_cout),
		.sum(u_comp_l0_p1_col19_sum));
	FullAdder u_comp_l0_p1_col20 (
		.a(u_comp_l0_p1_col20_a),
		.b(u_comp_l0_p1_col20_b),
		.cin(u_comp_l0_p1_col20_cin),
		.cout(u_comp_l0_p1_col20_cout),
		.sum(u_comp_l0_p1_col20_sum));
	FullAdder u_comp_l0_p1_col21 (
		.a(u_comp_l0_p1_col21_a),
		.b(u_comp_l0_p1_col21_b),
		.cin(u_comp_l0_p1_col21_cin),
		.cout(u_comp_l0_p1_col21_cout),
		.sum(u_comp_l0_p1_col21_sum));
	FullAdder u_comp_l0_p1_col22 (
		.a(u_comp_l0_p1_col22_a),
		.b(u_comp_l0_p1_col22_b),
		.cin(u_comp_l0_p1_col22_cin),
		.cout(u_comp_l0_p1_col22_cout),
		.sum(u_comp_l0_p1_col22_sum));
	FullAdder u_comp_l0_p1_col23 (
		.a(u_comp_l0_p1_col23_a),
		.b(u_comp_l0_p1_col23_b),
		.cin(u_comp_l0_p1_col23_cin),
		.cout(u_comp_l0_p1_col23_cout),
		.sum(u_comp_l0_p1_col23_sum));
	FullAdder u_comp_l0_p1_col24 (
		.a(u_comp_l0_p1_col24_a),
		.b(u_comp_l0_p1_col24_b),
		.cin(u_comp_l0_p1_col24_cin),
		.cout(u_comp_l0_p1_col24_cout),
		.sum(u_comp_l0_p1_col24_sum));
	FullAdder u_comp_l0_p1_col25 (
		.a(u_comp_l0_p1_col25_a),
		.b(u_comp_l0_p1_col25_b),
		.cin(u_comp_l0_p1_col25_cin),
		.cout(u_comp_l0_p1_col25_cout),
		.sum(u_comp_l0_p1_col25_sum));
	FullAdder u_comp_l0_p1_col26 (
		.a(u_comp_l0_p1_col26_a),
		.b(u_comp_l0_p1_col26_b),
		.cin(u_comp_l0_p1_col26_cin),
		.cout(u_comp_l0_p1_col26_cout),
		.sum(u_comp_l0_p1_col26_sum));
	FullAdder u_comp_l0_p1_col27 (
		.a(u_comp_l0_p1_col27_a),
		.b(u_comp_l0_p1_col27_b),
		.cin(u_comp_l0_p1_col27_cin),
		.cout(u_comp_l0_p1_col27_cout),
		.sum(u_comp_l0_p1_col27_sum));
	FullAdder u_comp_l0_p1_col28 (
		.a(u_comp_l0_p1_col28_a),
		.b(u_comp_l0_p1_col28_b),
		.cin(u_comp_l0_p1_col28_cin),
		.cout(u_comp_l0_p1_col28_cout),
		.sum(u_comp_l0_p1_col28_sum));
	FullAdder u_comp_l0_p1_col29 (
		.a(u_comp_l0_p1_col29_a),
		.b(u_comp_l0_p1_col29_b),
		.cin(u_comp_l0_p1_col29_cin),
		.cout(u_comp_l0_p1_col29_cout),
		.sum(u_comp_l0_p1_col29_sum));
	FullAdder u_comp_l0_p1_col30 (
		.a(u_comp_l0_p1_col30_a),
		.b(u_comp_l0_p1_col30_b),
		.cin(u_comp_l0_p1_col30_cin),
		.cout(u_comp_l0_p1_col30_cout),
		.sum(u_comp_l0_p1_col30_sum));
	FullAdder u_comp_l0_p1_col31 (
		.a(u_comp_l0_p1_col31_a),
		.b(u_comp_l0_p1_col31_b),
		.cin(u_comp_l0_p1_col31_cin),
		.cout(comp_l0_p1_col31_cout),
		.sum(u_comp_l0_p1_col31_sum));
	FullAdder u_comp_l0_p2_col0 (
		.a(u_comp_l0_p2_col0_a),
		.b(u_comp_l0_p2_col0_b),
		.cin(u_comp_l0_p2_col0_cin),
		.cout(u_comp_l0_p2_col0_cout),
		.sum(u_comp_l0_p2_col0_sum));
	FullAdder u_comp_l0_p2_col1 (
		.a(u_comp_l0_p2_col1_a),
		.b(u_comp_l0_p2_col1_b),
		.cin(u_comp_l0_p2_col1_cin),
		.cout(u_comp_l0_p2_col1_cout),
		.sum(u_comp_l0_p2_col1_sum));
	FullAdder u_comp_l0_p2_col2 (
		.a(u_comp_l0_p2_col2_a),
		.b(u_comp_l0_p2_col2_b),
		.cin(u_comp_l0_p2_col2_cin),
		.cout(u_comp_l0_p2_col2_cout),
		.sum(u_comp_l0_p2_col2_sum));
	FullAdder u_comp_l0_p2_col3 (
		.a(u_comp_l0_p2_col3_a),
		.b(u_comp_l0_p2_col3_b),
		.cin(u_comp_l0_p2_col3_cin),
		.cout(u_comp_l0_p2_col3_cout),
		.sum(u_comp_l0_p2_col3_sum));
	FullAdder u_comp_l0_p2_col4 (
		.a(u_comp_l0_p2_col4_a),
		.b(u_comp_l0_p2_col4_b),
		.cin(u_comp_l0_p2_col4_cin),
		.cout(u_comp_l0_p2_col4_cout),
		.sum(u_comp_l0_p2_col4_sum));
	FullAdder u_comp_l0_p2_col5 (
		.a(u_comp_l0_p2_col5_a),
		.b(u_comp_l0_p2_col5_b),
		.cin(u_comp_l0_p2_col5_cin),
		.cout(u_comp_l0_p2_col5_cout),
		.sum(u_comp_l0_p2_col5_sum));
	FullAdder u_comp_l0_p2_col6 (
		.a(u_comp_l0_p2_col6_a),
		.b(u_comp_l0_p2_col6_b),
		.cin(u_comp_l0_p2_col6_cin),
		.cout(u_comp_l0_p2_col6_cout),
		.sum(u_comp_l0_p2_col6_sum));
	FullAdder u_comp_l0_p2_col7 (
		.a(u_comp_l0_p2_col7_a),
		.b(u_comp_l0_p2_col7_b),
		.cin(u_comp_l0_p2_col7_cin),
		.cout(u_comp_l0_p2_col7_cout),
		.sum(u_comp_l0_p2_col7_sum));
	FullAdder u_comp_l0_p2_col8 (
		.a(u_comp_l0_p2_col8_a),
		.b(u_comp_l0_p2_col8_b),
		.cin(u_comp_l0_p2_col8_cin),
		.cout(u_comp_l0_p2_col8_cout),
		.sum(u_comp_l0_p2_col8_sum));
	FullAdder u_comp_l0_p2_col9 (
		.a(u_comp_l0_p2_col9_a),
		.b(u_comp_l0_p2_col9_b),
		.cin(u_comp_l0_p2_col9_cin),
		.cout(u_comp_l0_p2_col9_cout),
		.sum(u_comp_l0_p2_col9_sum));
	FullAdder u_comp_l0_p2_col10 (
		.a(u_comp_l0_p2_col10_a),
		.b(u_comp_l0_p2_col10_b),
		.cin(u_comp_l0_p2_col10_cin),
		.cout(u_comp_l0_p2_col10_cout),
		.sum(u_comp_l0_p2_col10_sum));
	FullAdder u_comp_l0_p2_col11 (
		.a(u_comp_l0_p2_col11_a),
		.b(u_comp_l0_p2_col11_b),
		.cin(u_comp_l0_p2_col11_cin),
		.cout(u_comp_l0_p2_col11_cout),
		.sum(u_comp_l0_p2_col11_sum));
	FullAdder u_comp_l0_p2_col12 (
		.a(u_comp_l0_p2_col12_a),
		.b(u_comp_l0_p2_col12_b),
		.cin(u_comp_l0_p2_col12_cin),
		.cout(u_comp_l0_p2_col12_cout),
		.sum(u_comp_l0_p2_col12_sum));
	FullAdder u_comp_l0_p2_col13 (
		.a(u_comp_l0_p2_col13_a),
		.b(u_comp_l0_p2_col13_b),
		.cin(u_comp_l0_p2_col13_cin),
		.cout(u_comp_l0_p2_col13_cout),
		.sum(u_comp_l0_p2_col13_sum));
	FullAdder u_comp_l0_p2_col14 (
		.a(u_comp_l0_p2_col14_a),
		.b(u_comp_l0_p2_col14_b),
		.cin(u_comp_l0_p2_col14_cin),
		.cout(u_comp_l0_p2_col14_cout),
		.sum(u_comp_l0_p2_col14_sum));
	FullAdder u_comp_l0_p2_col15 (
		.a(u_comp_l0_p2_col15_a),
		.b(u_comp_l0_p2_col15_b),
		.cin(u_comp_l0_p2_col15_cin),
		.cout(u_comp_l0_p2_col15_cout),
		.sum(u_comp_l0_p2_col15_sum));
	FullAdder u_comp_l0_p2_col16 (
		.a(u_comp_l0_p2_col16_a),
		.b(u_comp_l0_p2_col16_b),
		.cin(u_comp_l0_p2_col16_cin),
		.cout(u_comp_l0_p2_col16_cout),
		.sum(u_comp_l0_p2_col16_sum));
	FullAdder u_comp_l0_p2_col17 (
		.a(u_comp_l0_p2_col17_a),
		.b(u_comp_l0_p2_col17_b),
		.cin(u_comp_l0_p2_col17_cin),
		.cout(u_comp_l0_p2_col17_cout),
		.sum(u_comp_l0_p2_col17_sum));
	FullAdder u_comp_l0_p2_col18 (
		.a(u_comp_l0_p2_col18_a),
		.b(u_comp_l0_p2_col18_b),
		.cin(u_comp_l0_p2_col18_cin),
		.cout(u_comp_l0_p2_col18_cout),
		.sum(u_comp_l0_p2_col18_sum));
	FullAdder u_comp_l0_p2_col19 (
		.a(u_comp_l0_p2_col19_a),
		.b(u_comp_l0_p2_col19_b),
		.cin(u_comp_l0_p2_col19_cin),
		.cout(u_comp_l0_p2_col19_cout),
		.sum(u_comp_l0_p2_col19_sum));
	FullAdder u_comp_l0_p2_col20 (
		.a(u_comp_l0_p2_col20_a),
		.b(u_comp_l0_p2_col20_b),
		.cin(u_comp_l0_p2_col20_cin),
		.cout(u_comp_l0_p2_col20_cout),
		.sum(u_comp_l0_p2_col20_sum));
	FullAdder u_comp_l0_p2_col21 (
		.a(u_comp_l0_p2_col21_a),
		.b(u_comp_l0_p2_col21_b),
		.cin(u_comp_l0_p2_col21_cin),
		.cout(u_comp_l0_p2_col21_cout),
		.sum(u_comp_l0_p2_col21_sum));
	FullAdder u_comp_l0_p2_col22 (
		.a(u_comp_l0_p2_col22_a),
		.b(u_comp_l0_p2_col22_b),
		.cin(u_comp_l0_p2_col22_cin),
		.cout(u_comp_l0_p2_col22_cout),
		.sum(u_comp_l0_p2_col22_sum));
	FullAdder u_comp_l0_p2_col23 (
		.a(u_comp_l0_p2_col23_a),
		.b(u_comp_l0_p2_col23_b),
		.cin(u_comp_l0_p2_col23_cin),
		.cout(u_comp_l0_p2_col23_cout),
		.sum(u_comp_l0_p2_col23_sum));
	FullAdder u_comp_l0_p2_col24 (
		.a(u_comp_l0_p2_col24_a),
		.b(u_comp_l0_p2_col24_b),
		.cin(u_comp_l0_p2_col24_cin),
		.cout(u_comp_l0_p2_col24_cout),
		.sum(u_comp_l0_p2_col24_sum));
	FullAdder u_comp_l0_p2_col25 (
		.a(u_comp_l0_p2_col25_a),
		.b(u_comp_l0_p2_col25_b),
		.cin(u_comp_l0_p2_col25_cin),
		.cout(u_comp_l0_p2_col25_cout),
		.sum(u_comp_l0_p2_col25_sum));
	FullAdder u_comp_l0_p2_col26 (
		.a(u_comp_l0_p2_col26_a),
		.b(u_comp_l0_p2_col26_b),
		.cin(u_comp_l0_p2_col26_cin),
		.cout(u_comp_l0_p2_col26_cout),
		.sum(u_comp_l0_p2_col26_sum));
	FullAdder u_comp_l0_p2_col27 (
		.a(u_comp_l0_p2_col27_a),
		.b(u_comp_l0_p2_col27_b),
		.cin(u_comp_l0_p2_col27_cin),
		.cout(u_comp_l0_p2_col27_cout),
		.sum(u_comp_l0_p2_col27_sum));
	FullAdder u_comp_l0_p2_col28 (
		.a(u_comp_l0_p2_col28_a),
		.b(u_comp_l0_p2_col28_b),
		.cin(u_comp_l0_p2_col28_cin),
		.cout(u_comp_l0_p2_col28_cout),
		.sum(u_comp_l0_p2_col28_sum));
	FullAdder u_comp_l0_p2_col29 (
		.a(u_comp_l0_p2_col29_a),
		.b(u_comp_l0_p2_col29_b),
		.cin(u_comp_l0_p2_col29_cin),
		.cout(u_comp_l0_p2_col29_cout),
		.sum(u_comp_l0_p2_col29_sum));
	FullAdder u_comp_l0_p2_col30 (
		.a(u_comp_l0_p2_col30_a),
		.b(u_comp_l0_p2_col30_b),
		.cin(u_comp_l0_p2_col30_cin),
		.cout(u_comp_l0_p2_col30_cout),
		.sum(u_comp_l0_p2_col30_sum));
	FullAdder u_comp_l0_p2_col31 (
		.a(u_comp_l0_p2_col31_a),
		.b(u_comp_l0_p2_col31_b),
		.cin(u_comp_l0_p2_col31_cin),
		.cout(comp_l0_p2_col31_cout),
		.sum(u_comp_l0_p2_col31_sum));
	FullAdder u_comp_l1_p0_col0 (
		.a(u_comp_l1_p0_col0_a),
		.b(u_comp_l1_p0_col0_b),
		.cin(u_comp_l1_p0_col0_cin),
		.cout(u_comp_l1_p0_col0_cout),
		.sum(u_comp_l1_p0_col0_sum));
	FullAdder u_comp_l1_p0_col1 (
		.a(u_comp_l1_p0_col1_a),
		.b(u_comp_l1_p0_col1_b),
		.cin(u_comp_l1_p0_col1_cin),
		.cout(u_comp_l1_p0_col1_cout),
		.sum(u_comp_l1_p0_col1_sum));
	FullAdder u_comp_l1_p0_col2 (
		.a(u_comp_l1_p0_col2_a),
		.b(u_comp_l1_p0_col2_b),
		.cin(u_comp_l1_p0_col2_cin),
		.cout(u_comp_l1_p0_col2_cout),
		.sum(u_comp_l1_p0_col2_sum));
	FullAdder u_comp_l1_p0_col3 (
		.a(u_comp_l1_p0_col3_a),
		.b(u_comp_l1_p0_col3_b),
		.cin(u_comp_l1_p0_col3_cin),
		.cout(u_comp_l1_p0_col3_cout),
		.sum(u_comp_l1_p0_col3_sum));
	FullAdder u_comp_l1_p0_col4 (
		.a(u_comp_l1_p0_col4_a),
		.b(u_comp_l1_p0_col4_b),
		.cin(u_comp_l1_p0_col4_cin),
		.cout(u_comp_l1_p0_col4_cout),
		.sum(u_comp_l1_p0_col4_sum));
	FullAdder u_comp_l1_p0_col5 (
		.a(u_comp_l1_p0_col5_a),
		.b(u_comp_l1_p0_col5_b),
		.cin(u_comp_l1_p0_col5_cin),
		.cout(u_comp_l1_p0_col5_cout),
		.sum(u_comp_l1_p0_col5_sum));
	FullAdder u_comp_l1_p0_col6 (
		.a(u_comp_l1_p0_col6_a),
		.b(u_comp_l1_p0_col6_b),
		.cin(u_comp_l1_p0_col6_cin),
		.cout(u_comp_l1_p0_col6_cout),
		.sum(u_comp_l1_p0_col6_sum));
	FullAdder u_comp_l1_p0_col7 (
		.a(u_comp_l1_p0_col7_a),
		.b(u_comp_l1_p0_col7_b),
		.cin(u_comp_l1_p0_col7_cin),
		.cout(u_comp_l1_p0_col7_cout),
		.sum(u_comp_l1_p0_col7_sum));
	FullAdder u_comp_l1_p0_col8 (
		.a(u_comp_l1_p0_col8_a),
		.b(u_comp_l1_p0_col8_b),
		.cin(u_comp_l1_p0_col8_cin),
		.cout(u_comp_l1_p0_col8_cout),
		.sum(u_comp_l1_p0_col8_sum));
	FullAdder u_comp_l1_p0_col9 (
		.a(u_comp_l1_p0_col9_a),
		.b(u_comp_l1_p0_col9_b),
		.cin(u_comp_l1_p0_col9_cin),
		.cout(u_comp_l1_p0_col9_cout),
		.sum(u_comp_l1_p0_col9_sum));
	FullAdder u_comp_l1_p0_col10 (
		.a(u_comp_l1_p0_col10_a),
		.b(u_comp_l1_p0_col10_b),
		.cin(u_comp_l1_p0_col10_cin),
		.cout(u_comp_l1_p0_col10_cout),
		.sum(u_comp_l1_p0_col10_sum));
	FullAdder u_comp_l1_p0_col11 (
		.a(u_comp_l1_p0_col11_a),
		.b(u_comp_l1_p0_col11_b),
		.cin(u_comp_l1_p0_col11_cin),
		.cout(u_comp_l1_p0_col11_cout),
		.sum(u_comp_l1_p0_col11_sum));
	FullAdder u_comp_l1_p0_col12 (
		.a(u_comp_l1_p0_col12_a),
		.b(u_comp_l1_p0_col12_b),
		.cin(u_comp_l1_p0_col12_cin),
		.cout(u_comp_l1_p0_col12_cout),
		.sum(u_comp_l1_p0_col12_sum));
	FullAdder u_comp_l1_p0_col13 (
		.a(u_comp_l1_p0_col13_a),
		.b(u_comp_l1_p0_col13_b),
		.cin(u_comp_l1_p0_col13_cin),
		.cout(u_comp_l1_p0_col13_cout),
		.sum(u_comp_l1_p0_col13_sum));
	FullAdder u_comp_l1_p0_col14 (
		.a(u_comp_l1_p0_col14_a),
		.b(u_comp_l1_p0_col14_b),
		.cin(u_comp_l1_p0_col14_cin),
		.cout(u_comp_l1_p0_col14_cout),
		.sum(u_comp_l1_p0_col14_sum));
	FullAdder u_comp_l1_p0_col15 (
		.a(u_comp_l1_p0_col15_a),
		.b(u_comp_l1_p0_col15_b),
		.cin(u_comp_l1_p0_col15_cin),
		.cout(u_comp_l1_p0_col15_cout),
		.sum(u_comp_l1_p0_col15_sum));
	FullAdder u_comp_l1_p0_col16 (
		.a(u_comp_l1_p0_col16_a),
		.b(u_comp_l1_p0_col16_b),
		.cin(u_comp_l1_p0_col16_cin),
		.cout(u_comp_l1_p0_col16_cout),
		.sum(u_comp_l1_p0_col16_sum));
	FullAdder u_comp_l1_p0_col17 (
		.a(u_comp_l1_p0_col17_a),
		.b(u_comp_l1_p0_col17_b),
		.cin(u_comp_l1_p0_col17_cin),
		.cout(u_comp_l1_p0_col17_cout),
		.sum(u_comp_l1_p0_col17_sum));
	FullAdder u_comp_l1_p0_col18 (
		.a(u_comp_l1_p0_col18_a),
		.b(u_comp_l1_p0_col18_b),
		.cin(u_comp_l1_p0_col18_cin),
		.cout(u_comp_l1_p0_col18_cout),
		.sum(u_comp_l1_p0_col18_sum));
	FullAdder u_comp_l1_p0_col19 (
		.a(u_comp_l1_p0_col19_a),
		.b(u_comp_l1_p0_col19_b),
		.cin(u_comp_l1_p0_col19_cin),
		.cout(u_comp_l1_p0_col19_cout),
		.sum(u_comp_l1_p0_col19_sum));
	FullAdder u_comp_l1_p0_col20 (
		.a(u_comp_l1_p0_col20_a),
		.b(u_comp_l1_p0_col20_b),
		.cin(u_comp_l1_p0_col20_cin),
		.cout(u_comp_l1_p0_col20_cout),
		.sum(u_comp_l1_p0_col20_sum));
	FullAdder u_comp_l1_p0_col21 (
		.a(u_comp_l1_p0_col21_a),
		.b(u_comp_l1_p0_col21_b),
		.cin(u_comp_l1_p0_col21_cin),
		.cout(u_comp_l1_p0_col21_cout),
		.sum(u_comp_l1_p0_col21_sum));
	FullAdder u_comp_l1_p0_col22 (
		.a(u_comp_l1_p0_col22_a),
		.b(u_comp_l1_p0_col22_b),
		.cin(u_comp_l1_p0_col22_cin),
		.cout(u_comp_l1_p0_col22_cout),
		.sum(u_comp_l1_p0_col22_sum));
	FullAdder u_comp_l1_p0_col23 (
		.a(u_comp_l1_p0_col23_a),
		.b(u_comp_l1_p0_col23_b),
		.cin(u_comp_l1_p0_col23_cin),
		.cout(u_comp_l1_p0_col23_cout),
		.sum(u_comp_l1_p0_col23_sum));
	FullAdder u_comp_l1_p0_col24 (
		.a(u_comp_l1_p0_col24_a),
		.b(u_comp_l1_p0_col24_b),
		.cin(u_comp_l1_p0_col24_cin),
		.cout(u_comp_l1_p0_col24_cout),
		.sum(u_comp_l1_p0_col24_sum));
	FullAdder u_comp_l1_p0_col25 (
		.a(u_comp_l1_p0_col25_a),
		.b(u_comp_l1_p0_col25_b),
		.cin(u_comp_l1_p0_col25_cin),
		.cout(u_comp_l1_p0_col25_cout),
		.sum(u_comp_l1_p0_col25_sum));
	FullAdder u_comp_l1_p0_col26 (
		.a(u_comp_l1_p0_col26_a),
		.b(u_comp_l1_p0_col26_b),
		.cin(u_comp_l1_p0_col26_cin),
		.cout(u_comp_l1_p0_col26_cout),
		.sum(u_comp_l1_p0_col26_sum));
	FullAdder u_comp_l1_p0_col27 (
		.a(u_comp_l1_p0_col27_a),
		.b(u_comp_l1_p0_col27_b),
		.cin(u_comp_l1_p0_col27_cin),
		.cout(u_comp_l1_p0_col27_cout),
		.sum(u_comp_l1_p0_col27_sum));
	FullAdder u_comp_l1_p0_col28 (
		.a(u_comp_l1_p0_col28_a),
		.b(u_comp_l1_p0_col28_b),
		.cin(u_comp_l1_p0_col28_cin),
		.cout(u_comp_l1_p0_col28_cout),
		.sum(u_comp_l1_p0_col28_sum));
	FullAdder u_comp_l1_p0_col29 (
		.a(u_comp_l1_p0_col29_a),
		.b(u_comp_l1_p0_col29_b),
		.cin(u_comp_l1_p0_col29_cin),
		.cout(u_comp_l1_p0_col29_cout),
		.sum(u_comp_l1_p0_col29_sum));
	FullAdder u_comp_l1_p0_col30 (
		.a(u_comp_l1_p0_col30_a),
		.b(u_comp_l1_p0_col30_b),
		.cin(u_comp_l1_p0_col30_cin),
		.cout(u_comp_l1_p0_col30_cout),
		.sum(u_comp_l1_p0_col30_sum));
	FullAdder u_comp_l1_p0_col31 (
		.a(u_comp_l1_p0_col31_a),
		.b(u_comp_l1_p0_col31_b),
		.cin(u_comp_l1_p0_col31_cin),
		.cout(comp_l1_p0_col31_cout),
		.sum(u_comp_l1_p0_col31_sum));
	FullAdder u_comp_l1_p1_col0 (
		.a(u_comp_l1_p1_col0_a),
		.b(u_comp_l1_p1_col0_b),
		.cin(u_comp_l1_p1_col0_cin),
		.cout(u_comp_l1_p1_col0_cout),
		.sum(u_comp_l1_p1_col0_sum));
	FullAdder u_comp_l1_p1_col1 (
		.a(u_comp_l1_p1_col1_a),
		.b(u_comp_l1_p1_col1_b),
		.cin(u_comp_l1_p1_col1_cin),
		.cout(u_comp_l1_p1_col1_cout),
		.sum(u_comp_l1_p1_col1_sum));
	FullAdder u_comp_l1_p1_col2 (
		.a(u_comp_l1_p1_col2_a),
		.b(u_comp_l1_p1_col2_b),
		.cin(u_comp_l1_p1_col2_cin),
		.cout(u_comp_l1_p1_col2_cout),
		.sum(u_comp_l1_p1_col2_sum));
	FullAdder u_comp_l1_p1_col3 (
		.a(u_comp_l1_p1_col3_a),
		.b(u_comp_l1_p1_col3_b),
		.cin(u_comp_l1_p1_col3_cin),
		.cout(u_comp_l1_p1_col3_cout),
		.sum(u_comp_l1_p1_col3_sum));
	FullAdder u_comp_l1_p1_col4 (
		.a(u_comp_l1_p1_col4_a),
		.b(u_comp_l1_p1_col4_b),
		.cin(u_comp_l1_p1_col4_cin),
		.cout(u_comp_l1_p1_col4_cout),
		.sum(u_comp_l1_p1_col4_sum));
	FullAdder u_comp_l1_p1_col5 (
		.a(u_comp_l1_p1_col5_a),
		.b(u_comp_l1_p1_col5_b),
		.cin(u_comp_l1_p1_col5_cin),
		.cout(u_comp_l1_p1_col5_cout),
		.sum(u_comp_l1_p1_col5_sum));
	FullAdder u_comp_l1_p1_col6 (
		.a(u_comp_l1_p1_col6_a),
		.b(u_comp_l1_p1_col6_b),
		.cin(u_comp_l1_p1_col6_cin),
		.cout(u_comp_l1_p1_col6_cout),
		.sum(u_comp_l1_p1_col6_sum));
	FullAdder u_comp_l1_p1_col7 (
		.a(u_comp_l1_p1_col7_a),
		.b(u_comp_l1_p1_col7_b),
		.cin(u_comp_l1_p1_col7_cin),
		.cout(u_comp_l1_p1_col7_cout),
		.sum(u_comp_l1_p1_col7_sum));
	FullAdder u_comp_l1_p1_col8 (
		.a(u_comp_l1_p1_col8_a),
		.b(u_comp_l1_p1_col8_b),
		.cin(u_comp_l1_p1_col8_cin),
		.cout(u_comp_l1_p1_col8_cout),
		.sum(u_comp_l1_p1_col8_sum));
	FullAdder u_comp_l1_p1_col9 (
		.a(u_comp_l1_p1_col9_a),
		.b(u_comp_l1_p1_col9_b),
		.cin(u_comp_l1_p1_col9_cin),
		.cout(u_comp_l1_p1_col9_cout),
		.sum(u_comp_l1_p1_col9_sum));
	FullAdder u_comp_l1_p1_col10 (
		.a(u_comp_l1_p1_col10_a),
		.b(u_comp_l1_p1_col10_b),
		.cin(u_comp_l1_p1_col10_cin),
		.cout(u_comp_l1_p1_col10_cout),
		.sum(u_comp_l1_p1_col10_sum));
	FullAdder u_comp_l1_p1_col11 (
		.a(u_comp_l1_p1_col11_a),
		.b(u_comp_l1_p1_col11_b),
		.cin(u_comp_l1_p1_col11_cin),
		.cout(u_comp_l1_p1_col11_cout),
		.sum(u_comp_l1_p1_col11_sum));
	FullAdder u_comp_l1_p1_col12 (
		.a(u_comp_l1_p1_col12_a),
		.b(u_comp_l1_p1_col12_b),
		.cin(u_comp_l1_p1_col12_cin),
		.cout(u_comp_l1_p1_col12_cout),
		.sum(u_comp_l1_p1_col12_sum));
	FullAdder u_comp_l1_p1_col13 (
		.a(u_comp_l1_p1_col13_a),
		.b(u_comp_l1_p1_col13_b),
		.cin(u_comp_l1_p1_col13_cin),
		.cout(u_comp_l1_p1_col13_cout),
		.sum(u_comp_l1_p1_col13_sum));
	FullAdder u_comp_l1_p1_col14 (
		.a(u_comp_l1_p1_col14_a),
		.b(u_comp_l1_p1_col14_b),
		.cin(u_comp_l1_p1_col14_cin),
		.cout(u_comp_l1_p1_col14_cout),
		.sum(u_comp_l1_p1_col14_sum));
	FullAdder u_comp_l1_p1_col15 (
		.a(u_comp_l1_p1_col15_a),
		.b(u_comp_l1_p1_col15_b),
		.cin(u_comp_l1_p1_col15_cin),
		.cout(u_comp_l1_p1_col15_cout),
		.sum(u_comp_l1_p1_col15_sum));
	FullAdder u_comp_l1_p1_col16 (
		.a(u_comp_l1_p1_col16_a),
		.b(u_comp_l1_p1_col16_b),
		.cin(u_comp_l1_p1_col16_cin),
		.cout(u_comp_l1_p1_col16_cout),
		.sum(u_comp_l1_p1_col16_sum));
	FullAdder u_comp_l1_p1_col17 (
		.a(u_comp_l1_p1_col17_a),
		.b(u_comp_l1_p1_col17_b),
		.cin(u_comp_l1_p1_col17_cin),
		.cout(u_comp_l1_p1_col17_cout),
		.sum(u_comp_l1_p1_col17_sum));
	FullAdder u_comp_l1_p1_col18 (
		.a(u_comp_l1_p1_col18_a),
		.b(u_comp_l1_p1_col18_b),
		.cin(u_comp_l1_p1_col18_cin),
		.cout(u_comp_l1_p1_col18_cout),
		.sum(u_comp_l1_p1_col18_sum));
	FullAdder u_comp_l1_p1_col19 (
		.a(u_comp_l1_p1_col19_a),
		.b(u_comp_l1_p1_col19_b),
		.cin(u_comp_l1_p1_col19_cin),
		.cout(u_comp_l1_p1_col19_cout),
		.sum(u_comp_l1_p1_col19_sum));
	FullAdder u_comp_l1_p1_col20 (
		.a(u_comp_l1_p1_col20_a),
		.b(u_comp_l1_p1_col20_b),
		.cin(u_comp_l1_p1_col20_cin),
		.cout(u_comp_l1_p1_col20_cout),
		.sum(u_comp_l1_p1_col20_sum));
	FullAdder u_comp_l1_p1_col21 (
		.a(u_comp_l1_p1_col21_a),
		.b(u_comp_l1_p1_col21_b),
		.cin(u_comp_l1_p1_col21_cin),
		.cout(u_comp_l1_p1_col21_cout),
		.sum(u_comp_l1_p1_col21_sum));
	FullAdder u_comp_l1_p1_col22 (
		.a(u_comp_l1_p1_col22_a),
		.b(u_comp_l1_p1_col22_b),
		.cin(u_comp_l1_p1_col22_cin),
		.cout(u_comp_l1_p1_col22_cout),
		.sum(u_comp_l1_p1_col22_sum));
	FullAdder u_comp_l1_p1_col23 (
		.a(u_comp_l1_p1_col23_a),
		.b(u_comp_l1_p1_col23_b),
		.cin(u_comp_l1_p1_col23_cin),
		.cout(u_comp_l1_p1_col23_cout),
		.sum(u_comp_l1_p1_col23_sum));
	FullAdder u_comp_l1_p1_col24 (
		.a(u_comp_l1_p1_col24_a),
		.b(u_comp_l1_p1_col24_b),
		.cin(u_comp_l1_p1_col24_cin),
		.cout(u_comp_l1_p1_col24_cout),
		.sum(u_comp_l1_p1_col24_sum));
	FullAdder u_comp_l1_p1_col25 (
		.a(u_comp_l1_p1_col25_a),
		.b(u_comp_l1_p1_col25_b),
		.cin(u_comp_l1_p1_col25_cin),
		.cout(u_comp_l1_p1_col25_cout),
		.sum(u_comp_l1_p1_col25_sum));
	FullAdder u_comp_l1_p1_col26 (
		.a(u_comp_l1_p1_col26_a),
		.b(u_comp_l1_p1_col26_b),
		.cin(u_comp_l1_p1_col26_cin),
		.cout(u_comp_l1_p1_col26_cout),
		.sum(u_comp_l1_p1_col26_sum));
	FullAdder u_comp_l1_p1_col27 (
		.a(u_comp_l1_p1_col27_a),
		.b(u_comp_l1_p1_col27_b),
		.cin(u_comp_l1_p1_col27_cin),
		.cout(u_comp_l1_p1_col27_cout),
		.sum(u_comp_l1_p1_col27_sum));
	FullAdder u_comp_l1_p1_col28 (
		.a(u_comp_l1_p1_col28_a),
		.b(u_comp_l1_p1_col28_b),
		.cin(u_comp_l1_p1_col28_cin),
		.cout(u_comp_l1_p1_col28_cout),
		.sum(u_comp_l1_p1_col28_sum));
	FullAdder u_comp_l1_p1_col29 (
		.a(u_comp_l1_p1_col29_a),
		.b(u_comp_l1_p1_col29_b),
		.cin(u_comp_l1_p1_col29_cin),
		.cout(u_comp_l1_p1_col29_cout),
		.sum(u_comp_l1_p1_col29_sum));
	FullAdder u_comp_l1_p1_col30 (
		.a(u_comp_l1_p1_col30_a),
		.b(u_comp_l1_p1_col30_b),
		.cin(u_comp_l1_p1_col30_cin),
		.cout(u_comp_l1_p1_col30_cout),
		.sum(u_comp_l1_p1_col30_sum));
	FullAdder u_comp_l1_p1_col31 (
		.a(u_comp_l1_p1_col31_a),
		.b(u_comp_l1_p1_col31_b),
		.cin(u_comp_l1_p1_col31_cin),
		.cout(comp_l1_p1_col31_cout),
		.sum(u_comp_l1_p1_col31_sum));
	FullAdder u_comp_l2_p0_col0 (
		.a(u_comp_l2_p0_col0_a),
		.b(u_comp_l2_p0_col0_b),
		.cin(u_comp_l2_p0_col0_cin),
		.cout(u_comp_l2_p0_col0_cout),
		.sum(u_comp_l2_p0_col0_sum));
	FullAdder u_comp_l2_p0_col1 (
		.a(u_comp_l2_p0_col1_a),
		.b(u_comp_l2_p0_col1_b),
		.cin(u_comp_l2_p0_col1_cin),
		.cout(u_comp_l2_p0_col1_cout),
		.sum(u_comp_l2_p0_col1_sum));
	FullAdder u_comp_l2_p0_col2 (
		.a(u_comp_l2_p0_col2_a),
		.b(u_comp_l2_p0_col2_b),
		.cin(u_comp_l2_p0_col2_cin),
		.cout(u_comp_l2_p0_col2_cout),
		.sum(u_comp_l2_p0_col2_sum));
	FullAdder u_comp_l2_p0_col3 (
		.a(u_comp_l2_p0_col3_a),
		.b(u_comp_l2_p0_col3_b),
		.cin(u_comp_l2_p0_col3_cin),
		.cout(u_comp_l2_p0_col3_cout),
		.sum(u_comp_l2_p0_col3_sum));
	FullAdder u_comp_l2_p0_col4 (
		.a(u_comp_l2_p0_col4_a),
		.b(u_comp_l2_p0_col4_b),
		.cin(u_comp_l2_p0_col4_cin),
		.cout(u_comp_l2_p0_col4_cout),
		.sum(u_comp_l2_p0_col4_sum));
	FullAdder u_comp_l2_p0_col5 (
		.a(u_comp_l2_p0_col5_a),
		.b(u_comp_l2_p0_col5_b),
		.cin(u_comp_l2_p0_col5_cin),
		.cout(u_comp_l2_p0_col5_cout),
		.sum(u_comp_l2_p0_col5_sum));
	FullAdder u_comp_l2_p0_col6 (
		.a(u_comp_l2_p0_col6_a),
		.b(u_comp_l2_p0_col6_b),
		.cin(u_comp_l2_p0_col6_cin),
		.cout(u_comp_l2_p0_col6_cout),
		.sum(u_comp_l2_p0_col6_sum));
	FullAdder u_comp_l2_p0_col7 (
		.a(u_comp_l2_p0_col7_a),
		.b(u_comp_l2_p0_col7_b),
		.cin(u_comp_l2_p0_col7_cin),
		.cout(u_comp_l2_p0_col7_cout),
		.sum(u_comp_l2_p0_col7_sum));
	FullAdder u_comp_l2_p0_col8 (
		.a(u_comp_l2_p0_col8_a),
		.b(u_comp_l2_p0_col8_b),
		.cin(u_comp_l2_p0_col8_cin),
		.cout(u_comp_l2_p0_col8_cout),
		.sum(u_comp_l2_p0_col8_sum));
	FullAdder u_comp_l2_p0_col9 (
		.a(u_comp_l2_p0_col9_a),
		.b(u_comp_l2_p0_col9_b),
		.cin(u_comp_l2_p0_col9_cin),
		.cout(u_comp_l2_p0_col9_cout),
		.sum(u_comp_l2_p0_col9_sum));
	FullAdder u_comp_l2_p0_col10 (
		.a(u_comp_l2_p0_col10_a),
		.b(u_comp_l2_p0_col10_b),
		.cin(u_comp_l2_p0_col10_cin),
		.cout(u_comp_l2_p0_col10_cout),
		.sum(u_comp_l2_p0_col10_sum));
	FullAdder u_comp_l2_p0_col11 (
		.a(u_comp_l2_p0_col11_a),
		.b(u_comp_l2_p0_col11_b),
		.cin(u_comp_l2_p0_col11_cin),
		.cout(u_comp_l2_p0_col11_cout),
		.sum(u_comp_l2_p0_col11_sum));
	FullAdder u_comp_l2_p0_col12 (
		.a(u_comp_l2_p0_col12_a),
		.b(u_comp_l2_p0_col12_b),
		.cin(u_comp_l2_p0_col12_cin),
		.cout(u_comp_l2_p0_col12_cout),
		.sum(u_comp_l2_p0_col12_sum));
	FullAdder u_comp_l2_p0_col13 (
		.a(u_comp_l2_p0_col13_a),
		.b(u_comp_l2_p0_col13_b),
		.cin(u_comp_l2_p0_col13_cin),
		.cout(u_comp_l2_p0_col13_cout),
		.sum(u_comp_l2_p0_col13_sum));
	FullAdder u_comp_l2_p0_col14 (
		.a(u_comp_l2_p0_col14_a),
		.b(u_comp_l2_p0_col14_b),
		.cin(u_comp_l2_p0_col14_cin),
		.cout(u_comp_l2_p0_col14_cout),
		.sum(u_comp_l2_p0_col14_sum));
	FullAdder u_comp_l2_p0_col15 (
		.a(u_comp_l2_p0_col15_a),
		.b(u_comp_l2_p0_col15_b),
		.cin(u_comp_l2_p0_col15_cin),
		.cout(u_comp_l2_p0_col15_cout),
		.sum(u_comp_l2_p0_col15_sum));
	FullAdder u_comp_l2_p0_col16 (
		.a(u_comp_l2_p0_col16_a),
		.b(u_comp_l2_p0_col16_b),
		.cin(u_comp_l2_p0_col16_cin),
		.cout(u_comp_l2_p0_col16_cout),
		.sum(u_comp_l2_p0_col16_sum));
	FullAdder u_comp_l2_p0_col17 (
		.a(u_comp_l2_p0_col17_a),
		.b(u_comp_l2_p0_col17_b),
		.cin(u_comp_l2_p0_col17_cin),
		.cout(u_comp_l2_p0_col17_cout),
		.sum(u_comp_l2_p0_col17_sum));
	FullAdder u_comp_l2_p0_col18 (
		.a(u_comp_l2_p0_col18_a),
		.b(u_comp_l2_p0_col18_b),
		.cin(u_comp_l2_p0_col18_cin),
		.cout(u_comp_l2_p0_col18_cout),
		.sum(u_comp_l2_p0_col18_sum));
	FullAdder u_comp_l2_p0_col19 (
		.a(u_comp_l2_p0_col19_a),
		.b(u_comp_l2_p0_col19_b),
		.cin(u_comp_l2_p0_col19_cin),
		.cout(u_comp_l2_p0_col19_cout),
		.sum(u_comp_l2_p0_col19_sum));
	FullAdder u_comp_l2_p0_col20 (
		.a(u_comp_l2_p0_col20_a),
		.b(u_comp_l2_p0_col20_b),
		.cin(u_comp_l2_p0_col20_cin),
		.cout(u_comp_l2_p0_col20_cout),
		.sum(u_comp_l2_p0_col20_sum));
	FullAdder u_comp_l2_p0_col21 (
		.a(u_comp_l2_p0_col21_a),
		.b(u_comp_l2_p0_col21_b),
		.cin(u_comp_l2_p0_col21_cin),
		.cout(u_comp_l2_p0_col21_cout),
		.sum(u_comp_l2_p0_col21_sum));
	FullAdder u_comp_l2_p0_col22 (
		.a(u_comp_l2_p0_col22_a),
		.b(u_comp_l2_p0_col22_b),
		.cin(u_comp_l2_p0_col22_cin),
		.cout(u_comp_l2_p0_col22_cout),
		.sum(u_comp_l2_p0_col22_sum));
	FullAdder u_comp_l2_p0_col23 (
		.a(u_comp_l2_p0_col23_a),
		.b(u_comp_l2_p0_col23_b),
		.cin(u_comp_l2_p0_col23_cin),
		.cout(u_comp_l2_p0_col23_cout),
		.sum(u_comp_l2_p0_col23_sum));
	FullAdder u_comp_l2_p0_col24 (
		.a(u_comp_l2_p0_col24_a),
		.b(u_comp_l2_p0_col24_b),
		.cin(u_comp_l2_p0_col24_cin),
		.cout(u_comp_l2_p0_col24_cout),
		.sum(u_comp_l2_p0_col24_sum));
	FullAdder u_comp_l2_p0_col25 (
		.a(u_comp_l2_p0_col25_a),
		.b(u_comp_l2_p0_col25_b),
		.cin(u_comp_l2_p0_col25_cin),
		.cout(u_comp_l2_p0_col25_cout),
		.sum(u_comp_l2_p0_col25_sum));
	FullAdder u_comp_l2_p0_col26 (
		.a(u_comp_l2_p0_col26_a),
		.b(u_comp_l2_p0_col26_b),
		.cin(u_comp_l2_p0_col26_cin),
		.cout(u_comp_l2_p0_col26_cout),
		.sum(u_comp_l2_p0_col26_sum));
	FullAdder u_comp_l2_p0_col27 (
		.a(u_comp_l2_p0_col27_a),
		.b(u_comp_l2_p0_col27_b),
		.cin(u_comp_l2_p0_col27_cin),
		.cout(u_comp_l2_p0_col27_cout),
		.sum(u_comp_l2_p0_col27_sum));
	FullAdder u_comp_l2_p0_col28 (
		.a(u_comp_l2_p0_col28_a),
		.b(u_comp_l2_p0_col28_b),
		.cin(u_comp_l2_p0_col28_cin),
		.cout(u_comp_l2_p0_col28_cout),
		.sum(u_comp_l2_p0_col28_sum));
	FullAdder u_comp_l2_p0_col29 (
		.a(u_comp_l2_p0_col29_a),
		.b(u_comp_l2_p0_col29_b),
		.cin(u_comp_l2_p0_col29_cin),
		.cout(u_comp_l2_p0_col29_cout),
		.sum(u_comp_l2_p0_col29_sum));
	FullAdder u_comp_l2_p0_col30 (
		.a(u_comp_l2_p0_col30_a),
		.b(u_comp_l2_p0_col30_b),
		.cin(u_comp_l2_p0_col30_cin),
		.cout(u_comp_l2_p0_col30_cout),
		.sum(u_comp_l2_p0_col30_sum));
	FullAdder u_comp_l2_p0_col31 (
		.a(u_comp_l2_p0_col31_a),
		.b(u_comp_l2_p0_col31_b),
		.cin(u_comp_l2_p0_col31_cin),
		.cout(comp_l2_p0_col31_cout),
		.sum(u_comp_l2_p0_col31_sum));
	FullAdder u_comp_l3_p0_col0 (
		.a(u_comp_l3_p0_col0_a),
		.b(u_comp_l3_p0_col0_b),
		.cin(u_comp_l3_p0_col0_cin),
		.cout(u_comp_l3_p0_col0_cout),
		.sum(u_comp_l3_p0_col0_sum));
	FullAdder u_comp_l3_p0_col1 (
		.a(u_comp_l3_p0_col1_a),
		.b(u_comp_l3_p0_col1_b),
		.cin(u_comp_l3_p0_col1_cin),
		.cout(u_comp_l3_p0_col1_cout),
		.sum(u_comp_l3_p0_col1_sum));
	FullAdder u_comp_l3_p0_col2 (
		.a(u_comp_l3_p0_col2_a),
		.b(u_comp_l3_p0_col2_b),
		.cin(u_comp_l3_p0_col2_cin),
		.cout(u_comp_l3_p0_col2_cout),
		.sum(u_comp_l3_p0_col2_sum));
	FullAdder u_comp_l3_p0_col3 (
		.a(u_comp_l3_p0_col3_a),
		.b(u_comp_l3_p0_col3_b),
		.cin(u_comp_l3_p0_col3_cin),
		.cout(u_comp_l3_p0_col3_cout),
		.sum(u_comp_l3_p0_col3_sum));
	FullAdder u_comp_l3_p0_col4 (
		.a(u_comp_l3_p0_col4_a),
		.b(u_comp_l3_p0_col4_b),
		.cin(u_comp_l3_p0_col4_cin),
		.cout(u_comp_l3_p0_col4_cout),
		.sum(u_comp_l3_p0_col4_sum));
	FullAdder u_comp_l3_p0_col5 (
		.a(u_comp_l3_p0_col5_a),
		.b(u_comp_l3_p0_col5_b),
		.cin(u_comp_l3_p0_col5_cin),
		.cout(u_comp_l3_p0_col5_cout),
		.sum(u_comp_l3_p0_col5_sum));
	FullAdder u_comp_l3_p0_col6 (
		.a(u_comp_l3_p0_col6_a),
		.b(u_comp_l3_p0_col6_b),
		.cin(u_comp_l3_p0_col6_cin),
		.cout(u_comp_l3_p0_col6_cout),
		.sum(u_comp_l3_p0_col6_sum));
	FullAdder u_comp_l3_p0_col7 (
		.a(u_comp_l3_p0_col7_a),
		.b(u_comp_l3_p0_col7_b),
		.cin(u_comp_l3_p0_col7_cin),
		.cout(u_comp_l3_p0_col7_cout),
		.sum(u_comp_l3_p0_col7_sum));
	FullAdder u_comp_l3_p0_col8 (
		.a(u_comp_l3_p0_col8_a),
		.b(u_comp_l3_p0_col8_b),
		.cin(u_comp_l3_p0_col8_cin),
		.cout(u_comp_l3_p0_col8_cout),
		.sum(u_comp_l3_p0_col8_sum));
	FullAdder u_comp_l3_p0_col9 (
		.a(u_comp_l3_p0_col9_a),
		.b(u_comp_l3_p0_col9_b),
		.cin(u_comp_l3_p0_col9_cin),
		.cout(u_comp_l3_p0_col9_cout),
		.sum(u_comp_l3_p0_col9_sum));
	FullAdder u_comp_l3_p0_col10 (
		.a(u_comp_l3_p0_col10_a),
		.b(u_comp_l3_p0_col10_b),
		.cin(u_comp_l3_p0_col10_cin),
		.cout(u_comp_l3_p0_col10_cout),
		.sum(u_comp_l3_p0_col10_sum));
	FullAdder u_comp_l3_p0_col11 (
		.a(u_comp_l3_p0_col11_a),
		.b(u_comp_l3_p0_col11_b),
		.cin(u_comp_l3_p0_col11_cin),
		.cout(u_comp_l3_p0_col11_cout),
		.sum(u_comp_l3_p0_col11_sum));
	FullAdder u_comp_l3_p0_col12 (
		.a(u_comp_l3_p0_col12_a),
		.b(u_comp_l3_p0_col12_b),
		.cin(u_comp_l3_p0_col12_cin),
		.cout(u_comp_l3_p0_col12_cout),
		.sum(u_comp_l3_p0_col12_sum));
	FullAdder u_comp_l3_p0_col13 (
		.a(u_comp_l3_p0_col13_a),
		.b(u_comp_l3_p0_col13_b),
		.cin(u_comp_l3_p0_col13_cin),
		.cout(u_comp_l3_p0_col13_cout),
		.sum(u_comp_l3_p0_col13_sum));
	FullAdder u_comp_l3_p0_col14 (
		.a(u_comp_l3_p0_col14_a),
		.b(u_comp_l3_p0_col14_b),
		.cin(u_comp_l3_p0_col14_cin),
		.cout(u_comp_l3_p0_col14_cout),
		.sum(u_comp_l3_p0_col14_sum));
	FullAdder u_comp_l3_p0_col15 (
		.a(u_comp_l3_p0_col15_a),
		.b(u_comp_l3_p0_col15_b),
		.cin(u_comp_l3_p0_col15_cin),
		.cout(u_comp_l3_p0_col15_cout),
		.sum(u_comp_l3_p0_col15_sum));
	FullAdder u_comp_l3_p0_col16 (
		.a(u_comp_l3_p0_col16_a),
		.b(u_comp_l3_p0_col16_b),
		.cin(u_comp_l3_p0_col16_cin),
		.cout(u_comp_l3_p0_col16_cout),
		.sum(u_comp_l3_p0_col16_sum));
	FullAdder u_comp_l3_p0_col17 (
		.a(u_comp_l3_p0_col17_a),
		.b(u_comp_l3_p0_col17_b),
		.cin(u_comp_l3_p0_col17_cin),
		.cout(u_comp_l3_p0_col17_cout),
		.sum(u_comp_l3_p0_col17_sum));
	FullAdder u_comp_l3_p0_col18 (
		.a(u_comp_l3_p0_col18_a),
		.b(u_comp_l3_p0_col18_b),
		.cin(u_comp_l3_p0_col18_cin),
		.cout(u_comp_l3_p0_col18_cout),
		.sum(u_comp_l3_p0_col18_sum));
	FullAdder u_comp_l3_p0_col19 (
		.a(u_comp_l3_p0_col19_a),
		.b(u_comp_l3_p0_col19_b),
		.cin(u_comp_l3_p0_col19_cin),
		.cout(u_comp_l3_p0_col19_cout),
		.sum(u_comp_l3_p0_col19_sum));
	FullAdder u_comp_l3_p0_col20 (
		.a(u_comp_l3_p0_col20_a),
		.b(u_comp_l3_p0_col20_b),
		.cin(u_comp_l3_p0_col20_cin),
		.cout(u_comp_l3_p0_col20_cout),
		.sum(u_comp_l3_p0_col20_sum));
	FullAdder u_comp_l3_p0_col21 (
		.a(u_comp_l3_p0_col21_a),
		.b(u_comp_l3_p0_col21_b),
		.cin(u_comp_l3_p0_col21_cin),
		.cout(u_comp_l3_p0_col21_cout),
		.sum(u_comp_l3_p0_col21_sum));
	FullAdder u_comp_l3_p0_col22 (
		.a(u_comp_l3_p0_col22_a),
		.b(u_comp_l3_p0_col22_b),
		.cin(u_comp_l3_p0_col22_cin),
		.cout(u_comp_l3_p0_col22_cout),
		.sum(u_comp_l3_p0_col22_sum));
	FullAdder u_comp_l3_p0_col23 (
		.a(u_comp_l3_p0_col23_a),
		.b(u_comp_l3_p0_col23_b),
		.cin(u_comp_l3_p0_col23_cin),
		.cout(u_comp_l3_p0_col23_cout),
		.sum(u_comp_l3_p0_col23_sum));
	FullAdder u_comp_l3_p0_col24 (
		.a(u_comp_l3_p0_col24_a),
		.b(u_comp_l3_p0_col24_b),
		.cin(u_comp_l3_p0_col24_cin),
		.cout(u_comp_l3_p0_col24_cout),
		.sum(u_comp_l3_p0_col24_sum));
	FullAdder u_comp_l3_p0_col25 (
		.a(u_comp_l3_p0_col25_a),
		.b(u_comp_l3_p0_col25_b),
		.cin(u_comp_l3_p0_col25_cin),
		.cout(u_comp_l3_p0_col25_cout),
		.sum(u_comp_l3_p0_col25_sum));
	FullAdder u_comp_l3_p0_col26 (
		.a(u_comp_l3_p0_col26_a),
		.b(u_comp_l3_p0_col26_b),
		.cin(u_comp_l3_p0_col26_cin),
		.cout(u_comp_l3_p0_col26_cout),
		.sum(u_comp_l3_p0_col26_sum));
	FullAdder u_comp_l3_p0_col27 (
		.a(u_comp_l3_p0_col27_a),
		.b(u_comp_l3_p0_col27_b),
		.cin(u_comp_l3_p0_col27_cin),
		.cout(u_comp_l3_p0_col27_cout),
		.sum(u_comp_l3_p0_col27_sum));
	FullAdder u_comp_l3_p0_col28 (
		.a(u_comp_l3_p0_col28_a),
		.b(u_comp_l3_p0_col28_b),
		.cin(u_comp_l3_p0_col28_cin),
		.cout(u_comp_l3_p0_col28_cout),
		.sum(u_comp_l3_p0_col28_sum));
	FullAdder u_comp_l3_p0_col29 (
		.a(u_comp_l3_p0_col29_a),
		.b(u_comp_l3_p0_col29_b),
		.cin(u_comp_l3_p0_col29_cin),
		.cout(u_comp_l3_p0_col29_cout),
		.sum(u_comp_l3_p0_col29_sum));
	FullAdder u_comp_l3_p0_col30 (
		.a(u_comp_l3_p0_col30_a),
		.b(u_comp_l3_p0_col30_b),
		.cin(u_comp_l3_p0_col30_cin),
		.cout(u_comp_l3_p0_col30_cout),
		.sum(u_comp_l3_p0_col30_sum));
	FullAdder u_comp_l3_p0_col31 (
		.a(u_comp_l3_p0_col31_a),
		.b(u_comp_l3_p0_col31_b),
		.cin(u_comp_l3_p0_col31_cin),
		.cout(comp_l3_p0_col31_cout),
		.sum(u_comp_l3_p0_col31_sum));
	FullAdder u_comp_l4_p0_col0 (
		.a(u_comp_l4_p0_col0_a),
		.b(u_comp_l4_p0_col0_b),
		.cin(u_comp_l4_p0_col0_cin),
		.cout(u_comp_l4_p0_col0_cout),
		.sum(u_comp_l4_p0_col0_sum));
	FullAdder u_comp_l4_p0_col1 (
		.a(u_comp_l4_p0_col1_a),
		.b(u_comp_l4_p0_col1_b),
		.cin(u_comp_l4_p0_col1_cin),
		.cout(u_comp_l4_p0_col1_cout),
		.sum(u_comp_l4_p0_col1_sum));
	FullAdder u_comp_l4_p0_col2 (
		.a(u_comp_l4_p0_col2_a),
		.b(u_comp_l4_p0_col2_b),
		.cin(u_comp_l4_p0_col2_cin),
		.cout(u_comp_l4_p0_col2_cout),
		.sum(u_comp_l4_p0_col2_sum));
	FullAdder u_comp_l4_p0_col3 (
		.a(u_comp_l4_p0_col3_a),
		.b(u_comp_l4_p0_col3_b),
		.cin(u_comp_l4_p0_col3_cin),
		.cout(u_comp_l4_p0_col3_cout),
		.sum(u_comp_l4_p0_col3_sum));
	FullAdder u_comp_l4_p0_col4 (
		.a(u_comp_l4_p0_col4_a),
		.b(u_comp_l4_p0_col4_b),
		.cin(u_comp_l4_p0_col4_cin),
		.cout(u_comp_l4_p0_col4_cout),
		.sum(u_comp_l4_p0_col4_sum));
	FullAdder u_comp_l4_p0_col5 (
		.a(u_comp_l4_p0_col5_a),
		.b(u_comp_l4_p0_col5_b),
		.cin(u_comp_l4_p0_col5_cin),
		.cout(u_comp_l4_p0_col5_cout),
		.sum(u_comp_l4_p0_col5_sum));
	FullAdder u_comp_l4_p0_col6 (
		.a(u_comp_l4_p0_col6_a),
		.b(u_comp_l4_p0_col6_b),
		.cin(u_comp_l4_p0_col6_cin),
		.cout(u_comp_l4_p0_col6_cout),
		.sum(u_comp_l4_p0_col6_sum));
	FullAdder u_comp_l4_p0_col7 (
		.a(u_comp_l4_p0_col7_a),
		.b(u_comp_l4_p0_col7_b),
		.cin(u_comp_l4_p0_col7_cin),
		.cout(u_comp_l4_p0_col7_cout),
		.sum(u_comp_l4_p0_col7_sum));
	FullAdder u_comp_l4_p0_col8 (
		.a(u_comp_l4_p0_col8_a),
		.b(u_comp_l4_p0_col8_b),
		.cin(u_comp_l4_p0_col8_cin),
		.cout(u_comp_l4_p0_col8_cout),
		.sum(u_comp_l4_p0_col8_sum));
	FullAdder u_comp_l4_p0_col9 (
		.a(u_comp_l4_p0_col9_a),
		.b(u_comp_l4_p0_col9_b),
		.cin(u_comp_l4_p0_col9_cin),
		.cout(u_comp_l4_p0_col9_cout),
		.sum(u_comp_l4_p0_col9_sum));
	FullAdder u_comp_l4_p0_col10 (
		.a(u_comp_l4_p0_col10_a),
		.b(u_comp_l4_p0_col10_b),
		.cin(u_comp_l4_p0_col10_cin),
		.cout(u_comp_l4_p0_col10_cout),
		.sum(u_comp_l4_p0_col10_sum));
	FullAdder u_comp_l4_p0_col11 (
		.a(u_comp_l4_p0_col11_a),
		.b(u_comp_l4_p0_col11_b),
		.cin(u_comp_l4_p0_col11_cin),
		.cout(u_comp_l4_p0_col11_cout),
		.sum(u_comp_l4_p0_col11_sum));
	FullAdder u_comp_l4_p0_col12 (
		.a(u_comp_l4_p0_col12_a),
		.b(u_comp_l4_p0_col12_b),
		.cin(u_comp_l4_p0_col12_cin),
		.cout(u_comp_l4_p0_col12_cout),
		.sum(u_comp_l4_p0_col12_sum));
	FullAdder u_comp_l4_p0_col13 (
		.a(u_comp_l4_p0_col13_a),
		.b(u_comp_l4_p0_col13_b),
		.cin(u_comp_l4_p0_col13_cin),
		.cout(u_comp_l4_p0_col13_cout),
		.sum(u_comp_l4_p0_col13_sum));
	FullAdder u_comp_l4_p0_col14 (
		.a(u_comp_l4_p0_col14_a),
		.b(u_comp_l4_p0_col14_b),
		.cin(u_comp_l4_p0_col14_cin),
		.cout(u_comp_l4_p0_col14_cout),
		.sum(u_comp_l4_p0_col14_sum));
	FullAdder u_comp_l4_p0_col15 (
		.a(u_comp_l4_p0_col15_a),
		.b(u_comp_l4_p0_col15_b),
		.cin(u_comp_l4_p0_col15_cin),
		.cout(u_comp_l4_p0_col15_cout),
		.sum(u_comp_l4_p0_col15_sum));
	FullAdder u_comp_l4_p0_col16 (
		.a(u_comp_l4_p0_col16_a),
		.b(u_comp_l4_p0_col16_b),
		.cin(u_comp_l4_p0_col16_cin),
		.cout(u_comp_l4_p0_col16_cout),
		.sum(u_comp_l4_p0_col16_sum));
	FullAdder u_comp_l4_p0_col17 (
		.a(u_comp_l4_p0_col17_a),
		.b(u_comp_l4_p0_col17_b),
		.cin(u_comp_l4_p0_col17_cin),
		.cout(u_comp_l4_p0_col17_cout),
		.sum(u_comp_l4_p0_col17_sum));
	FullAdder u_comp_l4_p0_col18 (
		.a(u_comp_l4_p0_col18_a),
		.b(u_comp_l4_p0_col18_b),
		.cin(u_comp_l4_p0_col18_cin),
		.cout(u_comp_l4_p0_col18_cout),
		.sum(u_comp_l4_p0_col18_sum));
	FullAdder u_comp_l4_p0_col19 (
		.a(u_comp_l4_p0_col19_a),
		.b(u_comp_l4_p0_col19_b),
		.cin(u_comp_l4_p0_col19_cin),
		.cout(u_comp_l4_p0_col19_cout),
		.sum(u_comp_l4_p0_col19_sum));
	FullAdder u_comp_l4_p0_col20 (
		.a(u_comp_l4_p0_col20_a),
		.b(u_comp_l4_p0_col20_b),
		.cin(u_comp_l4_p0_col20_cin),
		.cout(u_comp_l4_p0_col20_cout),
		.sum(u_comp_l4_p0_col20_sum));
	FullAdder u_comp_l4_p0_col21 (
		.a(u_comp_l4_p0_col21_a),
		.b(u_comp_l4_p0_col21_b),
		.cin(u_comp_l4_p0_col21_cin),
		.cout(u_comp_l4_p0_col21_cout),
		.sum(u_comp_l4_p0_col21_sum));
	FullAdder u_comp_l4_p0_col22 (
		.a(u_comp_l4_p0_col22_a),
		.b(u_comp_l4_p0_col22_b),
		.cin(u_comp_l4_p0_col22_cin),
		.cout(u_comp_l4_p0_col22_cout),
		.sum(u_comp_l4_p0_col22_sum));
	FullAdder u_comp_l4_p0_col23 (
		.a(u_comp_l4_p0_col23_a),
		.b(u_comp_l4_p0_col23_b),
		.cin(u_comp_l4_p0_col23_cin),
		.cout(u_comp_l4_p0_col23_cout),
		.sum(u_comp_l4_p0_col23_sum));
	FullAdder u_comp_l4_p0_col24 (
		.a(u_comp_l4_p0_col24_a),
		.b(u_comp_l4_p0_col24_b),
		.cin(u_comp_l4_p0_col24_cin),
		.cout(u_comp_l4_p0_col24_cout),
		.sum(u_comp_l4_p0_col24_sum));
	FullAdder u_comp_l4_p0_col25 (
		.a(u_comp_l4_p0_col25_a),
		.b(u_comp_l4_p0_col25_b),
		.cin(u_comp_l4_p0_col25_cin),
		.cout(u_comp_l4_p0_col25_cout),
		.sum(u_comp_l4_p0_col25_sum));
	FullAdder u_comp_l4_p0_col26 (
		.a(u_comp_l4_p0_col26_a),
		.b(u_comp_l4_p0_col26_b),
		.cin(u_comp_l4_p0_col26_cin),
		.cout(u_comp_l4_p0_col26_cout),
		.sum(u_comp_l4_p0_col26_sum));
	FullAdder u_comp_l4_p0_col27 (
		.a(u_comp_l4_p0_col27_a),
		.b(u_comp_l4_p0_col27_b),
		.cin(u_comp_l4_p0_col27_cin),
		.cout(u_comp_l4_p0_col27_cout),
		.sum(u_comp_l4_p0_col27_sum));
	FullAdder u_comp_l4_p0_col28 (
		.a(u_comp_l4_p0_col28_a),
		.b(u_comp_l4_p0_col28_b),
		.cin(u_comp_l4_p0_col28_cin),
		.cout(u_comp_l4_p0_col28_cout),
		.sum(u_comp_l4_p0_col28_sum));
	FullAdder u_comp_l4_p0_col29 (
		.a(u_comp_l4_p0_col29_a),
		.b(u_comp_l4_p0_col29_b),
		.cin(u_comp_l4_p0_col29_cin),
		.cout(u_comp_l4_p0_col29_cout),
		.sum(u_comp_l4_p0_col29_sum));
	FullAdder u_comp_l4_p0_col30 (
		.a(u_comp_l4_p0_col30_a),
		.b(u_comp_l4_p0_col30_b),
		.cin(u_comp_l4_p0_col30_cin),
		.cout(u_comp_l4_p0_col30_cout),
		.sum(u_comp_l4_p0_col30_sum));
	FullAdder u_comp_l4_p0_col31 (
		.a(u_comp_l4_p0_col31_a),
		.b(u_comp_l4_p0_col31_b),
		.cin(u_comp_l4_p0_col31_cin),
		.cout(comp_l4_p0_col31_cout),
		.sum(u_comp_l4_p0_col31_sum));

endmodule
//[UHDL]Content End [md5:6e927582602471e237b52f7140ea2183]

